typedef logic [31:0] data_t;

module median_57_292_26 (
    input logic clk,
    input data_t data_0,
    input data_t data_1,
    input data_t data_2,
    input data_t data_3,
    input data_t data_4,
    input data_t data_5,
    input data_t data_6,
    input data_t data_7,
    input data_t data_8,
    input data_t data_9,
    input data_t data_10,
    input data_t data_11,
    input data_t data_12,
    input data_t data_13,
    input data_t data_14,
    input data_t data_15,
    input data_t data_16,
    input data_t data_17,
    input data_t data_18,
    input data_t data_19,
    input data_t data_20,
    input data_t data_21,
    input data_t data_22,
    input data_t data_23,
    input data_t data_24,
    input data_t data_25,
    input data_t data_26,
    input data_t data_27,
    input data_t data_28,
    input data_t data_29,
    input data_t data_30,
    input data_t data_31,
    input data_t data_32,
    input data_t data_33,
    input data_t data_34,
    input data_t data_35,
    input data_t data_36,
    input data_t data_37,
    input data_t data_38,
    input data_t data_39,
    input data_t data_40,
    input data_t data_41,
    input data_t data_42,
    input data_t data_43,
    input data_t data_44,
    input data_t data_45,
    input data_t data_46,
    input data_t data_47,
    input data_t data_48,
    input data_t data_49,
    input data_t data_50,
    input data_t data_51,
    input data_t data_52,
    input data_t data_53,
    input data_t data_54,
    input data_t data_55,
    input data_t data_56,
    output data_t sort_0,
    output data_t sort_1,
    output data_t sort_2,
    output data_t sort_3,
    output data_t sort_4,
    output data_t sort_5,
    output data_t sort_6,
    output data_t sort_7,
    output data_t sort_8,
    output data_t sort_9,
    output data_t sort_10,
    output data_t sort_11,
    output data_t sort_12,
    output data_t sort_13,
    output data_t sort_14,
    output data_t sort_15,
    output data_t sort_16,
    output data_t sort_17,
    output data_t sort_18,
    output data_t sort_19,
    output data_t sort_20,
    output data_t sort_21,
    output data_t sort_22,
    output data_t sort_23,
    output data_t sort_24,
    output data_t sort_25,
    output data_t sort_26,
    output data_t sort_27,
    output data_t sort_28,
    output data_t sort_29,
    output data_t sort_30,
    output data_t sort_31,
    output data_t sort_32,
    output data_t sort_33,
    output data_t sort_34,
    output data_t sort_35,
    output data_t sort_36,
    output data_t sort_37,
    output data_t sort_38,
    output data_t sort_39,
    output data_t sort_40,
    output data_t sort_41,
    output data_t sort_42,
    output data_t sort_43,
    output data_t sort_44,
    output data_t sort_45,
    output data_t sort_46,
    output data_t sort_47,
    output data_t sort_48,
    output data_t sort_49,
    output data_t sort_50,
    output data_t sort_51,
    output data_t sort_52,
    output data_t sort_53,
    output data_t sort_54,
    output data_t sort_55,
    output data_t sort_56
);

     logic [31:0] stage_0_out_0;
     logic [31:0] stage_0_out_1;
     logic [31:0] stage_0_out_2;
     logic [31:0] stage_0_out_3;
     logic [31:0] stage_0_out_4;
     logic [31:0] stage_0_out_5;
     logic [31:0] stage_0_out_6;
     logic [31:0] stage_0_out_7;
     logic [31:0] stage_0_out_8;
     logic [31:0] stage_0_out_9;
     logic [31:0] stage_0_out_10;
     logic [31:0] stage_0_out_11;
     logic [31:0] stage_0_out_12;
     logic [31:0] stage_0_out_13;
     logic [31:0] stage_0_out_14;
     logic [31:0] stage_0_out_15;
     logic [31:0] stage_0_out_16;
     logic [31:0] stage_0_out_17;
     logic [31:0] stage_0_out_18;
     logic [31:0] stage_0_out_19;
     logic [31:0] stage_0_out_20;
     logic [31:0] stage_0_out_21;
     logic [31:0] stage_0_out_22;
     logic [31:0] stage_0_out_23;
     logic [31:0] stage_0_out_24;
     logic [31:0] stage_0_out_25;
     logic [31:0] stage_0_out_26;
     logic [31:0] stage_0_out_27;
     logic [31:0] stage_0_out_28;
     logic [31:0] stage_0_out_29;
     logic [31:0] stage_0_out_30;
     logic [31:0] stage_0_out_31;
     logic [31:0] stage_0_out_32;
     logic [31:0] stage_0_out_33;
     logic [31:0] stage_0_out_34;
     logic [31:0] stage_0_out_35;
     logic [31:0] stage_0_out_36;
     logic [31:0] stage_0_out_37;
     logic [31:0] stage_0_out_38;
     logic [31:0] stage_0_out_39;
     logic [31:0] stage_0_out_40;
     logic [31:0] stage_0_out_41;
     logic [31:0] stage_0_out_42;
     logic [31:0] stage_0_out_43;
     logic [31:0] stage_0_out_44;
     logic [31:0] stage_0_out_45;
     logic [31:0] stage_0_out_46;
     logic [31:0] stage_0_out_47;
     logic [31:0] stage_0_out_48;
     logic [31:0] stage_0_out_49;
     logic [31:0] stage_0_out_50;
     logic [31:0] stage_0_out_51;
     logic [31:0] stage_0_out_52;
     logic [31:0] stage_0_out_53;
     logic [31:0] stage_0_out_54;
     logic [31:0] stage_0_out_55;
     logic [31:0] stage_0_out_56;
     logic [31:0] stage_1_out_0;
     logic [31:0] stage_1_out_1;
     logic [31:0] stage_1_out_2;
     logic [31:0] stage_1_out_3;
     logic [31:0] stage_1_out_4;
     logic [31:0] stage_1_out_5;
     logic [31:0] stage_1_out_6;
     logic [31:0] stage_1_out_7;
     logic [31:0] stage_1_out_8;
     logic [31:0] stage_1_out_9;
     logic [31:0] stage_1_out_10;
     logic [31:0] stage_1_out_11;
     logic [31:0] stage_1_out_12;
     logic [31:0] stage_1_out_13;
     logic [31:0] stage_1_out_14;
     logic [31:0] stage_1_out_15;
     logic [31:0] stage_1_out_16;
     logic [31:0] stage_1_out_17;
     logic [31:0] stage_1_out_18;
     logic [31:0] stage_1_out_19;
     logic [31:0] stage_1_out_20;
     logic [31:0] stage_1_out_21;
     logic [31:0] stage_1_out_22;
     logic [31:0] stage_1_out_23;
     logic [31:0] stage_1_out_24;
     logic [31:0] stage_1_out_25;
     logic [31:0] stage_1_out_26;
     logic [31:0] stage_1_out_27;
     logic [31:0] stage_1_out_28;
     logic [31:0] stage_1_out_29;
     logic [31:0] stage_1_out_30;
     logic [31:0] stage_1_out_31;
     logic [31:0] stage_1_out_32;
     logic [31:0] stage_1_out_33;
     logic [31:0] stage_1_out_34;
     logic [31:0] stage_1_out_35;
     logic [31:0] stage_1_out_36;
     logic [31:0] stage_1_out_37;
     logic [31:0] stage_1_out_38;
     logic [31:0] stage_1_out_39;
     logic [31:0] stage_1_out_40;
     logic [31:0] stage_1_out_41;
     logic [31:0] stage_1_out_42;
     logic [31:0] stage_1_out_43;
     logic [31:0] stage_1_out_44;
     logic [31:0] stage_1_out_45;
     logic [31:0] stage_1_out_46;
     logic [31:0] stage_1_out_47;
     logic [31:0] stage_1_out_48;
     logic [31:0] stage_1_out_49;
     logic [31:0] stage_1_out_50;
     logic [31:0] stage_1_out_51;
     logic [31:0] stage_1_out_52;
     logic [31:0] stage_1_out_53;
     logic [31:0] stage_1_out_54;
     logic [31:0] stage_1_out_55;
     logic [31:0] stage_1_out_56;
     logic [31:0] stage_2_out_0;
     logic [31:0] stage_2_out_1;
     logic [31:0] stage_2_out_2;
     logic [31:0] stage_2_out_3;
     logic [31:0] stage_2_out_4;
     logic [31:0] stage_2_out_5;
     logic [31:0] stage_2_out_6;
     logic [31:0] stage_2_out_7;
     logic [31:0] stage_2_out_8;
     logic [31:0] stage_2_out_9;
     logic [31:0] stage_2_out_10;
     logic [31:0] stage_2_out_11;
     logic [31:0] stage_2_out_12;
     logic [31:0] stage_2_out_13;
     logic [31:0] stage_2_out_14;
     logic [31:0] stage_2_out_15;
     logic [31:0] stage_2_out_16;
     logic [31:0] stage_2_out_17;
     logic [31:0] stage_2_out_18;
     logic [31:0] stage_2_out_19;
     logic [31:0] stage_2_out_20;
     logic [31:0] stage_2_out_21;
     logic [31:0] stage_2_out_22;
     logic [31:0] stage_2_out_23;
     logic [31:0] stage_2_out_24;
     logic [31:0] stage_2_out_25;
     logic [31:0] stage_2_out_26;
     logic [31:0] stage_2_out_27;
     logic [31:0] stage_2_out_28;
     logic [31:0] stage_2_out_29;
     logic [31:0] stage_2_out_30;
     logic [31:0] stage_2_out_31;
     logic [31:0] stage_2_out_32;
     logic [31:0] stage_2_out_33;
     logic [31:0] stage_2_out_34;
     logic [31:0] stage_2_out_35;
     logic [31:0] stage_2_out_36;
     logic [31:0] stage_2_out_37;
     logic [31:0] stage_2_out_38;
     logic [31:0] stage_2_out_39;
     logic [31:0] stage_2_out_40;
     logic [31:0] stage_2_out_41;
     logic [31:0] stage_2_out_42;
     logic [31:0] stage_2_out_43;
     logic [31:0] stage_2_out_44;
     logic [31:0] stage_2_out_45;
     logic [31:0] stage_2_out_46;
     logic [31:0] stage_2_out_47;
     logic [31:0] stage_2_out_48;
     logic [31:0] stage_2_out_49;
     logic [31:0] stage_2_out_50;
     logic [31:0] stage_2_out_51;
     logic [31:0] stage_2_out_52;
     logic [31:0] stage_2_out_53;
     logic [31:0] stage_2_out_54;
     logic [31:0] stage_2_out_55;
     logic [31:0] stage_2_out_56;
     logic [31:0] stage_3_out_0;
     logic [31:0] stage_3_out_1;
     logic [31:0] stage_3_out_2;
     logic [31:0] stage_3_out_3;
     logic [31:0] stage_3_out_4;
     logic [31:0] stage_3_out_5;
     logic [31:0] stage_3_out_6;
     logic [31:0] stage_3_out_7;
     logic [31:0] stage_3_out_8;
     logic [31:0] stage_3_out_9;
     logic [31:0] stage_3_out_10;
     logic [31:0] stage_3_out_11;
     logic [31:0] stage_3_out_12;
     logic [31:0] stage_3_out_13;
     logic [31:0] stage_3_out_14;
     logic [31:0] stage_3_out_15;
     logic [31:0] stage_3_out_16;
     logic [31:0] stage_3_out_17;
     logic [31:0] stage_3_out_18;
     logic [31:0] stage_3_out_19;
     logic [31:0] stage_3_out_20;
     logic [31:0] stage_3_out_21;
     logic [31:0] stage_3_out_22;
     logic [31:0] stage_3_out_23;
     logic [31:0] stage_3_out_24;
     logic [31:0] stage_3_out_25;
     logic [31:0] stage_3_out_26;
     logic [31:0] stage_3_out_27;
     logic [31:0] stage_3_out_28;
     logic [31:0] stage_3_out_29;
     logic [31:0] stage_3_out_30;
     logic [31:0] stage_3_out_31;
     logic [31:0] stage_3_out_32;
     logic [31:0] stage_3_out_33;
     logic [31:0] stage_3_out_34;
     logic [31:0] stage_3_out_35;
     logic [31:0] stage_3_out_36;
     logic [31:0] stage_3_out_37;
     logic [31:0] stage_3_out_38;
     logic [31:0] stage_3_out_39;
     logic [31:0] stage_3_out_40;
     logic [31:0] stage_3_out_41;
     logic [31:0] stage_3_out_42;
     logic [31:0] stage_3_out_43;
     logic [31:0] stage_3_out_44;
     logic [31:0] stage_3_out_45;
     logic [31:0] stage_3_out_46;
     logic [31:0] stage_3_out_47;
     logic [31:0] stage_3_out_48;
     logic [31:0] stage_3_out_49;
     logic [31:0] stage_3_out_50;
     logic [31:0] stage_3_out_51;
     logic [31:0] stage_3_out_52;
     logic [31:0] stage_3_out_53;
     logic [31:0] stage_3_out_54;
     logic [31:0] stage_3_out_55;
     logic [31:0] stage_3_out_56;
     logic [31:0] stage_4_out_0;
     logic [31:0] stage_4_out_1;
     logic [31:0] stage_4_out_2;
     logic [31:0] stage_4_out_3;
     logic [31:0] stage_4_out_4;
     logic [31:0] stage_4_out_5;
     logic [31:0] stage_4_out_6;
     logic [31:0] stage_4_out_7;
     logic [31:0] stage_4_out_8;
     logic [31:0] stage_4_out_9;
     logic [31:0] stage_4_out_10;
     logic [31:0] stage_4_out_11;
     logic [31:0] stage_4_out_12;
     logic [31:0] stage_4_out_13;
     logic [31:0] stage_4_out_14;
     logic [31:0] stage_4_out_15;
     logic [31:0] stage_4_out_16;
     logic [31:0] stage_4_out_17;
     logic [31:0] stage_4_out_18;
     logic [31:0] stage_4_out_19;
     logic [31:0] stage_4_out_20;
     logic [31:0] stage_4_out_21;
     logic [31:0] stage_4_out_22;
     logic [31:0] stage_4_out_23;
     logic [31:0] stage_4_out_24;
     logic [31:0] stage_4_out_25;
     logic [31:0] stage_4_out_26;
     logic [31:0] stage_4_out_27;
     logic [31:0] stage_4_out_28;
     logic [31:0] stage_4_out_29;
     logic [31:0] stage_4_out_30;
     logic [31:0] stage_4_out_31;
     logic [31:0] stage_4_out_32;
     logic [31:0] stage_4_out_33;
     logic [31:0] stage_4_out_34;
     logic [31:0] stage_4_out_35;
     logic [31:0] stage_4_out_36;
     logic [31:0] stage_4_out_37;
     logic [31:0] stage_4_out_38;
     logic [31:0] stage_4_out_39;
     logic [31:0] stage_4_out_40;
     logic [31:0] stage_4_out_41;
     logic [31:0] stage_4_out_42;
     logic [31:0] stage_4_out_43;
     logic [31:0] stage_4_out_44;
     logic [31:0] stage_4_out_45;
     logic [31:0] stage_4_out_46;
     logic [31:0] stage_4_out_47;
     logic [31:0] stage_4_out_48;
     logic [31:0] stage_4_out_49;
     logic [31:0] stage_4_out_50;
     logic [31:0] stage_4_out_51;
     logic [31:0] stage_4_out_52;
     logic [31:0] stage_4_out_53;
     logic [31:0] stage_4_out_54;
     logic [31:0] stage_4_out_55;
     logic [31:0] stage_4_out_56;
     logic [31:0] stage_5_out_0;
     logic [31:0] stage_5_out_1;
     logic [31:0] stage_5_out_2;
     logic [31:0] stage_5_out_3;
     logic [31:0] stage_5_out_4;
     logic [31:0] stage_5_out_5;
     logic [31:0] stage_5_out_6;
     logic [31:0] stage_5_out_7;
     logic [31:0] stage_5_out_8;
     logic [31:0] stage_5_out_9;
     logic [31:0] stage_5_out_10;
     logic [31:0] stage_5_out_11;
     logic [31:0] stage_5_out_12;
     logic [31:0] stage_5_out_13;
     logic [31:0] stage_5_out_14;
     logic [31:0] stage_5_out_15;
     logic [31:0] stage_5_out_16;
     logic [31:0] stage_5_out_17;
     logic [31:0] stage_5_out_18;
     logic [31:0] stage_5_out_19;
     logic [31:0] stage_5_out_20;
     logic [31:0] stage_5_out_21;
     logic [31:0] stage_5_out_22;
     logic [31:0] stage_5_out_23;
     logic [31:0] stage_5_out_24;
     logic [31:0] stage_5_out_25;
     logic [31:0] stage_5_out_26;
     logic [31:0] stage_5_out_27;
     logic [31:0] stage_5_out_28;
     logic [31:0] stage_5_out_29;
     logic [31:0] stage_5_out_30;
     logic [31:0] stage_5_out_31;
     logic [31:0] stage_5_out_32;
     logic [31:0] stage_5_out_33;
     logic [31:0] stage_5_out_34;
     logic [31:0] stage_5_out_35;
     logic [31:0] stage_5_out_36;
     logic [31:0] stage_5_out_37;
     logic [31:0] stage_5_out_38;
     logic [31:0] stage_5_out_39;
     logic [31:0] stage_5_out_40;
     logic [31:0] stage_5_out_41;
     logic [31:0] stage_5_out_42;
     logic [31:0] stage_5_out_43;
     logic [31:0] stage_5_out_44;
     logic [31:0] stage_5_out_45;
     logic [31:0] stage_5_out_46;
     logic [31:0] stage_5_out_47;
     logic [31:0] stage_5_out_48;
     logic [31:0] stage_5_out_49;
     logic [31:0] stage_5_out_50;
     logic [31:0] stage_5_out_51;
     logic [31:0] stage_5_out_52;
     logic [31:0] stage_5_out_53;
     logic [31:0] stage_5_out_54;
     logic [31:0] stage_5_out_55;
     logic [31:0] stage_5_out_56;
     logic [31:0] stage_6_out_0;
     logic [31:0] stage_6_out_1;
     logic [31:0] stage_6_out_2;
     logic [31:0] stage_6_out_3;
     logic [31:0] stage_6_out_4;
     logic [31:0] stage_6_out_5;
     logic [31:0] stage_6_out_6;
     logic [31:0] stage_6_out_7;
     logic [31:0] stage_6_out_8;
     logic [31:0] stage_6_out_9;
     logic [31:0] stage_6_out_10;
     logic [31:0] stage_6_out_11;
     logic [31:0] stage_6_out_12;
     logic [31:0] stage_6_out_13;
     logic [31:0] stage_6_out_14;
     logic [31:0] stage_6_out_15;
     logic [31:0] stage_6_out_16;
     logic [31:0] stage_6_out_17;
     logic [31:0] stage_6_out_18;
     logic [31:0] stage_6_out_19;
     logic [31:0] stage_6_out_20;
     logic [31:0] stage_6_out_21;
     logic [31:0] stage_6_out_22;
     logic [31:0] stage_6_out_23;
     logic [31:0] stage_6_out_24;
     logic [31:0] stage_6_out_25;
     logic [31:0] stage_6_out_26;
     logic [31:0] stage_6_out_27;
     logic [31:0] stage_6_out_28;
     logic [31:0] stage_6_out_29;
     logic [31:0] stage_6_out_30;
     logic [31:0] stage_6_out_31;
     logic [31:0] stage_6_out_32;
     logic [31:0] stage_6_out_33;
     logic [31:0] stage_6_out_34;
     logic [31:0] stage_6_out_35;
     logic [31:0] stage_6_out_36;
     logic [31:0] stage_6_out_37;
     logic [31:0] stage_6_out_38;
     logic [31:0] stage_6_out_39;
     logic [31:0] stage_6_out_40;
     logic [31:0] stage_6_out_41;
     logic [31:0] stage_6_out_42;
     logic [31:0] stage_6_out_43;
     logic [31:0] stage_6_out_44;
     logic [31:0] stage_6_out_45;
     logic [31:0] stage_6_out_46;
     logic [31:0] stage_6_out_47;
     logic [31:0] stage_6_out_48;
     logic [31:0] stage_6_out_49;
     logic [31:0] stage_6_out_50;
     logic [31:0] stage_6_out_51;
     logic [31:0] stage_6_out_52;
     logic [31:0] stage_6_out_53;
     logic [31:0] stage_6_out_54;
     logic [31:0] stage_6_out_55;
     logic [31:0] stage_6_out_56;
     logic [31:0] stage_7_out_0;
     logic [31:0] stage_7_out_1;
     logic [31:0] stage_7_out_2;
     logic [31:0] stage_7_out_3;
     logic [31:0] stage_7_out_4;
     logic [31:0] stage_7_out_5;
     logic [31:0] stage_7_out_6;
     logic [31:0] stage_7_out_7;
     logic [31:0] stage_7_out_8;
     logic [31:0] stage_7_out_9;
     logic [31:0] stage_7_out_10;
     logic [31:0] stage_7_out_11;
     logic [31:0] stage_7_out_12;
     logic [31:0] stage_7_out_13;
     logic [31:0] stage_7_out_14;
     logic [31:0] stage_7_out_15;
     logic [31:0] stage_7_out_16;
     logic [31:0] stage_7_out_17;
     logic [31:0] stage_7_out_18;
     logic [31:0] stage_7_out_19;
     logic [31:0] stage_7_out_20;
     logic [31:0] stage_7_out_21;
     logic [31:0] stage_7_out_22;
     logic [31:0] stage_7_out_23;
     logic [31:0] stage_7_out_24;
     logic [31:0] stage_7_out_25;
     logic [31:0] stage_7_out_26;
     logic [31:0] stage_7_out_27;
     logic [31:0] stage_7_out_28;
     logic [31:0] stage_7_out_29;
     logic [31:0] stage_7_out_30;
     logic [31:0] stage_7_out_31;
     logic [31:0] stage_7_out_32;
     logic [31:0] stage_7_out_33;
     logic [31:0] stage_7_out_34;
     logic [31:0] stage_7_out_35;
     logic [31:0] stage_7_out_36;
     logic [31:0] stage_7_out_37;
     logic [31:0] stage_7_out_38;
     logic [31:0] stage_7_out_39;
     logic [31:0] stage_7_out_40;
     logic [31:0] stage_7_out_41;
     logic [31:0] stage_7_out_42;
     logic [31:0] stage_7_out_43;
     logic [31:0] stage_7_out_44;
     logic [31:0] stage_7_out_45;
     logic [31:0] stage_7_out_46;
     logic [31:0] stage_7_out_47;
     logic [31:0] stage_7_out_48;
     logic [31:0] stage_7_out_49;
     logic [31:0] stage_7_out_50;
     logic [31:0] stage_7_out_51;
     logic [31:0] stage_7_out_52;
     logic [31:0] stage_7_out_53;
     logic [31:0] stage_7_out_54;
     logic [31:0] stage_7_out_55;
     logic [31:0] stage_7_out_56;
     logic [31:0] stage_8_out_0;
     logic [31:0] stage_8_out_1;
     logic [31:0] stage_8_out_2;
     logic [31:0] stage_8_out_3;
     logic [31:0] stage_8_out_4;
     logic [31:0] stage_8_out_5;
     logic [31:0] stage_8_out_6;
     logic [31:0] stage_8_out_7;
     logic [31:0] stage_8_out_8;
     logic [31:0] stage_8_out_9;
     logic [31:0] stage_8_out_10;
     logic [31:0] stage_8_out_11;
     logic [31:0] stage_8_out_12;
     logic [31:0] stage_8_out_13;
     logic [31:0] stage_8_out_14;
     logic [31:0] stage_8_out_15;
     logic [31:0] stage_8_out_16;
     logic [31:0] stage_8_out_17;
     logic [31:0] stage_8_out_18;
     logic [31:0] stage_8_out_19;
     logic [31:0] stage_8_out_20;
     logic [31:0] stage_8_out_21;
     logic [31:0] stage_8_out_22;
     logic [31:0] stage_8_out_23;
     logic [31:0] stage_8_out_24;
     logic [31:0] stage_8_out_25;
     logic [31:0] stage_8_out_26;
     logic [31:0] stage_8_out_27;
     logic [31:0] stage_8_out_28;
     logic [31:0] stage_8_out_29;
     logic [31:0] stage_8_out_30;
     logic [31:0] stage_8_out_31;
     logic [31:0] stage_8_out_32;
     logic [31:0] stage_8_out_33;
     logic [31:0] stage_8_out_34;
     logic [31:0] stage_8_out_35;
     logic [31:0] stage_8_out_36;
     logic [31:0] stage_8_out_37;
     logic [31:0] stage_8_out_38;
     logic [31:0] stage_8_out_39;
     logic [31:0] stage_8_out_40;
     logic [31:0] stage_8_out_41;
     logic [31:0] stage_8_out_42;
     logic [31:0] stage_8_out_43;
     logic [31:0] stage_8_out_44;
     logic [31:0] stage_8_out_45;
     logic [31:0] stage_8_out_46;
     logic [31:0] stage_8_out_47;
     logic [31:0] stage_8_out_48;
     logic [31:0] stage_8_out_49;
     logic [31:0] stage_8_out_50;
     logic [31:0] stage_8_out_51;
     logic [31:0] stage_8_out_52;
     logic [31:0] stage_8_out_53;
     logic [31:0] stage_8_out_54;
     logic [31:0] stage_8_out_55;
     logic [31:0] stage_8_out_56;
     logic [31:0] stage_9_out_0;
     logic [31:0] stage_9_out_1;
     logic [31:0] stage_9_out_2;
     logic [31:0] stage_9_out_3;
     logic [31:0] stage_9_out_4;
     logic [31:0] stage_9_out_5;
     logic [31:0] stage_9_out_6;
     logic [31:0] stage_9_out_7;
     logic [31:0] stage_9_out_8;
     logic [31:0] stage_9_out_9;
     logic [31:0] stage_9_out_10;
     logic [31:0] stage_9_out_11;
     logic [31:0] stage_9_out_12;
     logic [31:0] stage_9_out_13;
     logic [31:0] stage_9_out_14;
     logic [31:0] stage_9_out_15;
     logic [31:0] stage_9_out_16;
     logic [31:0] stage_9_out_17;
     logic [31:0] stage_9_out_18;
     logic [31:0] stage_9_out_19;
     logic [31:0] stage_9_out_20;
     logic [31:0] stage_9_out_21;
     logic [31:0] stage_9_out_22;
     logic [31:0] stage_9_out_23;
     logic [31:0] stage_9_out_24;
     logic [31:0] stage_9_out_25;
     logic [31:0] stage_9_out_26;
     logic [31:0] stage_9_out_27;
     logic [31:0] stage_9_out_28;
     logic [31:0] stage_9_out_29;
     logic [31:0] stage_9_out_30;
     logic [31:0] stage_9_out_31;
     logic [31:0] stage_9_out_32;
     logic [31:0] stage_9_out_33;
     logic [31:0] stage_9_out_34;
     logic [31:0] stage_9_out_35;
     logic [31:0] stage_9_out_36;
     logic [31:0] stage_9_out_37;
     logic [31:0] stage_9_out_38;
     logic [31:0] stage_9_out_39;
     logic [31:0] stage_9_out_40;
     logic [31:0] stage_9_out_41;
     logic [31:0] stage_9_out_42;
     logic [31:0] stage_9_out_43;
     logic [31:0] stage_9_out_44;
     logic [31:0] stage_9_out_45;
     logic [31:0] stage_9_out_46;
     logic [31:0] stage_9_out_47;
     logic [31:0] stage_9_out_48;
     logic [31:0] stage_9_out_49;
     logic [31:0] stage_9_out_50;
     logic [31:0] stage_9_out_51;
     logic [31:0] stage_9_out_52;
     logic [31:0] stage_9_out_53;
     logic [31:0] stage_9_out_54;
     logic [31:0] stage_9_out_55;
     logic [31:0] stage_9_out_56;
     logic [31:0] stage_10_out_0;
     logic [31:0] stage_10_out_1;
     logic [31:0] stage_10_out_2;
     logic [31:0] stage_10_out_3;
     logic [31:0] stage_10_out_4;
     logic [31:0] stage_10_out_5;
     logic [31:0] stage_10_out_6;
     logic [31:0] stage_10_out_7;
     logic [31:0] stage_10_out_8;
     logic [31:0] stage_10_out_9;
     logic [31:0] stage_10_out_10;
     logic [31:0] stage_10_out_11;
     logic [31:0] stage_10_out_12;
     logic [31:0] stage_10_out_13;
     logic [31:0] stage_10_out_14;
     logic [31:0] stage_10_out_15;
     logic [31:0] stage_10_out_16;
     logic [31:0] stage_10_out_17;
     logic [31:0] stage_10_out_18;
     logic [31:0] stage_10_out_19;
     logic [31:0] stage_10_out_20;
     logic [31:0] stage_10_out_21;
     logic [31:0] stage_10_out_22;
     logic [31:0] stage_10_out_23;
     logic [31:0] stage_10_out_24;
     logic [31:0] stage_10_out_25;
     logic [31:0] stage_10_out_26;
     logic [31:0] stage_10_out_27;
     logic [31:0] stage_10_out_28;
     logic [31:0] stage_10_out_29;
     logic [31:0] stage_10_out_30;
     logic [31:0] stage_10_out_31;
     logic [31:0] stage_10_out_32;
     logic [31:0] stage_10_out_33;
     logic [31:0] stage_10_out_34;
     logic [31:0] stage_10_out_35;
     logic [31:0] stage_10_out_36;
     logic [31:0] stage_10_out_37;
     logic [31:0] stage_10_out_38;
     logic [31:0] stage_10_out_39;
     logic [31:0] stage_10_out_40;
     logic [31:0] stage_10_out_41;
     logic [31:0] stage_10_out_42;
     logic [31:0] stage_10_out_43;
     logic [31:0] stage_10_out_44;
     logic [31:0] stage_10_out_45;
     logic [31:0] stage_10_out_46;
     logic [31:0] stage_10_out_47;
     logic [31:0] stage_10_out_48;
     logic [31:0] stage_10_out_49;
     logic [31:0] stage_10_out_50;
     logic [31:0] stage_10_out_51;
     logic [31:0] stage_10_out_52;
     logic [31:0] stage_10_out_53;
     logic [31:0] stage_10_out_54;
     logic [31:0] stage_10_out_55;
     logic [31:0] stage_10_out_56;
     logic [31:0] stage_11_out_0;
     logic [31:0] stage_11_out_1;
     logic [31:0] stage_11_out_2;
     logic [31:0] stage_11_out_3;
     logic [31:0] stage_11_out_4;
     logic [31:0] stage_11_out_5;
     logic [31:0] stage_11_out_6;
     logic [31:0] stage_11_out_7;
     logic [31:0] stage_11_out_8;
     logic [31:0] stage_11_out_9;
     logic [31:0] stage_11_out_10;
     logic [31:0] stage_11_out_11;
     logic [31:0] stage_11_out_12;
     logic [31:0] stage_11_out_13;
     logic [31:0] stage_11_out_14;
     logic [31:0] stage_11_out_15;
     logic [31:0] stage_11_out_16;
     logic [31:0] stage_11_out_17;
     logic [31:0] stage_11_out_18;
     logic [31:0] stage_11_out_19;
     logic [31:0] stage_11_out_20;
     logic [31:0] stage_11_out_21;
     logic [31:0] stage_11_out_22;
     logic [31:0] stage_11_out_23;
     logic [31:0] stage_11_out_24;
     logic [31:0] stage_11_out_25;
     logic [31:0] stage_11_out_26;
     logic [31:0] stage_11_out_27;
     logic [31:0] stage_11_out_28;
     logic [31:0] stage_11_out_29;
     logic [31:0] stage_11_out_30;
     logic [31:0] stage_11_out_31;
     logic [31:0] stage_11_out_32;
     logic [31:0] stage_11_out_33;
     logic [31:0] stage_11_out_34;
     logic [31:0] stage_11_out_35;
     logic [31:0] stage_11_out_36;
     logic [31:0] stage_11_out_37;
     logic [31:0] stage_11_out_38;
     logic [31:0] stage_11_out_39;
     logic [31:0] stage_11_out_40;
     logic [31:0] stage_11_out_41;
     logic [31:0] stage_11_out_42;
     logic [31:0] stage_11_out_43;
     logic [31:0] stage_11_out_44;
     logic [31:0] stage_11_out_45;
     logic [31:0] stage_11_out_46;
     logic [31:0] stage_11_out_47;
     logic [31:0] stage_11_out_48;
     logic [31:0] stage_11_out_49;
     logic [31:0] stage_11_out_50;
     logic [31:0] stage_11_out_51;
     logic [31:0] stage_11_out_52;
     logic [31:0] stage_11_out_53;
     logic [31:0] stage_11_out_54;
     logic [31:0] stage_11_out_55;
     logic [31:0] stage_11_out_56;
     logic [31:0] stage_12_out_0;
     logic [31:0] stage_12_out_1;
     logic [31:0] stage_12_out_2;
     logic [31:0] stage_12_out_3;
     logic [31:0] stage_12_out_4;
     logic [31:0] stage_12_out_5;
     logic [31:0] stage_12_out_6;
     logic [31:0] stage_12_out_7;
     logic [31:0] stage_12_out_8;
     logic [31:0] stage_12_out_9;
     logic [31:0] stage_12_out_10;
     logic [31:0] stage_12_out_11;
     logic [31:0] stage_12_out_12;
     logic [31:0] stage_12_out_13;
     logic [31:0] stage_12_out_14;
     logic [31:0] stage_12_out_15;
     logic [31:0] stage_12_out_16;
     logic [31:0] stage_12_out_17;
     logic [31:0] stage_12_out_18;
     logic [31:0] stage_12_out_19;
     logic [31:0] stage_12_out_20;
     logic [31:0] stage_12_out_21;
     logic [31:0] stage_12_out_22;
     logic [31:0] stage_12_out_23;
     logic [31:0] stage_12_out_24;
     logic [31:0] stage_12_out_25;
     logic [31:0] stage_12_out_26;
     logic [31:0] stage_12_out_27;
     logic [31:0] stage_12_out_28;
     logic [31:0] stage_12_out_29;
     logic [31:0] stage_12_out_30;
     logic [31:0] stage_12_out_31;
     logic [31:0] stage_12_out_32;
     logic [31:0] stage_12_out_33;
     logic [31:0] stage_12_out_34;
     logic [31:0] stage_12_out_35;
     logic [31:0] stage_12_out_36;
     logic [31:0] stage_12_out_37;
     logic [31:0] stage_12_out_38;
     logic [31:0] stage_12_out_39;
     logic [31:0] stage_12_out_40;
     logic [31:0] stage_12_out_41;
     logic [31:0] stage_12_out_42;
     logic [31:0] stage_12_out_43;
     logic [31:0] stage_12_out_44;
     logic [31:0] stage_12_out_45;
     logic [31:0] stage_12_out_46;
     logic [31:0] stage_12_out_47;
     logic [31:0] stage_12_out_48;
     logic [31:0] stage_12_out_49;
     logic [31:0] stage_12_out_50;
     logic [31:0] stage_12_out_51;
     logic [31:0] stage_12_out_52;
     logic [31:0] stage_12_out_53;
     logic [31:0] stage_12_out_54;
     logic [31:0] stage_12_out_55;
     logic [31:0] stage_12_out_56;
     logic [31:0] stage_13_out_0;
     logic [31:0] stage_13_out_1;
     logic [31:0] stage_13_out_2;
     logic [31:0] stage_13_out_3;
     logic [31:0] stage_13_out_4;
     logic [31:0] stage_13_out_5;
     logic [31:0] stage_13_out_6;
     logic [31:0] stage_13_out_7;
     logic [31:0] stage_13_out_8;
     logic [31:0] stage_13_out_9;
     logic [31:0] stage_13_out_10;
     logic [31:0] stage_13_out_11;
     logic [31:0] stage_13_out_12;
     logic [31:0] stage_13_out_13;
     logic [31:0] stage_13_out_14;
     logic [31:0] stage_13_out_15;
     logic [31:0] stage_13_out_16;
     logic [31:0] stage_13_out_17;
     logic [31:0] stage_13_out_18;
     logic [31:0] stage_13_out_19;
     logic [31:0] stage_13_out_20;
     logic [31:0] stage_13_out_21;
     logic [31:0] stage_13_out_22;
     logic [31:0] stage_13_out_23;
     logic [31:0] stage_13_out_24;
     logic [31:0] stage_13_out_25;
     logic [31:0] stage_13_out_26;
     logic [31:0] stage_13_out_27;
     logic [31:0] stage_13_out_28;
     logic [31:0] stage_13_out_29;
     logic [31:0] stage_13_out_30;
     logic [31:0] stage_13_out_31;
     logic [31:0] stage_13_out_32;
     logic [31:0] stage_13_out_33;
     logic [31:0] stage_13_out_34;
     logic [31:0] stage_13_out_35;
     logic [31:0] stage_13_out_36;
     logic [31:0] stage_13_out_37;
     logic [31:0] stage_13_out_38;
     logic [31:0] stage_13_out_39;
     logic [31:0] stage_13_out_40;
     logic [31:0] stage_13_out_41;
     logic [31:0] stage_13_out_42;
     logic [31:0] stage_13_out_43;
     logic [31:0] stage_13_out_44;
     logic [31:0] stage_13_out_45;
     logic [31:0] stage_13_out_46;
     logic [31:0] stage_13_out_47;
     logic [31:0] stage_13_out_48;
     logic [31:0] stage_13_out_49;
     logic [31:0] stage_13_out_50;
     logic [31:0] stage_13_out_51;
     logic [31:0] stage_13_out_52;
     logic [31:0] stage_13_out_53;
     logic [31:0] stage_13_out_54;
     logic [31:0] stage_13_out_55;
     logic [31:0] stage_13_out_56;
     logic [31:0] stage_14_out_0;
     logic [31:0] stage_14_out_1;
     logic [31:0] stage_14_out_2;
     logic [31:0] stage_14_out_3;
     logic [31:0] stage_14_out_4;
     logic [31:0] stage_14_out_5;
     logic [31:0] stage_14_out_6;
     logic [31:0] stage_14_out_7;
     logic [31:0] stage_14_out_8;
     logic [31:0] stage_14_out_9;
     logic [31:0] stage_14_out_10;
     logic [31:0] stage_14_out_11;
     logic [31:0] stage_14_out_12;
     logic [31:0] stage_14_out_13;
     logic [31:0] stage_14_out_14;
     logic [31:0] stage_14_out_15;
     logic [31:0] stage_14_out_16;
     logic [31:0] stage_14_out_17;
     logic [31:0] stage_14_out_18;
     logic [31:0] stage_14_out_19;
     logic [31:0] stage_14_out_20;
     logic [31:0] stage_14_out_21;
     logic [31:0] stage_14_out_22;
     logic [31:0] stage_14_out_23;
     logic [31:0] stage_14_out_24;
     logic [31:0] stage_14_out_25;
     logic [31:0] stage_14_out_26;
     logic [31:0] stage_14_out_27;
     logic [31:0] stage_14_out_28;
     logic [31:0] stage_14_out_29;
     logic [31:0] stage_14_out_30;
     logic [31:0] stage_14_out_31;
     logic [31:0] stage_14_out_32;
     logic [31:0] stage_14_out_33;
     logic [31:0] stage_14_out_34;
     logic [31:0] stage_14_out_35;
     logic [31:0] stage_14_out_36;
     logic [31:0] stage_14_out_37;
     logic [31:0] stage_14_out_38;
     logic [31:0] stage_14_out_39;
     logic [31:0] stage_14_out_40;
     logic [31:0] stage_14_out_41;
     logic [31:0] stage_14_out_42;
     logic [31:0] stage_14_out_43;
     logic [31:0] stage_14_out_44;
     logic [31:0] stage_14_out_45;
     logic [31:0] stage_14_out_46;
     logic [31:0] stage_14_out_47;
     logic [31:0] stage_14_out_48;
     logic [31:0] stage_14_out_49;
     logic [31:0] stage_14_out_50;
     logic [31:0] stage_14_out_51;
     logic [31:0] stage_14_out_52;
     logic [31:0] stage_14_out_53;
     logic [31:0] stage_14_out_54;
     logic [31:0] stage_14_out_55;
     logic [31:0] stage_14_out_56;
     logic [31:0] stage_15_out_0;
     logic [31:0] stage_15_out_1;
     logic [31:0] stage_15_out_2;
     logic [31:0] stage_15_out_3;
     logic [31:0] stage_15_out_4;
     logic [31:0] stage_15_out_5;
     logic [31:0] stage_15_out_6;
     logic [31:0] stage_15_out_7;
     logic [31:0] stage_15_out_8;
     logic [31:0] stage_15_out_9;
     logic [31:0] stage_15_out_10;
     logic [31:0] stage_15_out_11;
     logic [31:0] stage_15_out_12;
     logic [31:0] stage_15_out_13;
     logic [31:0] stage_15_out_14;
     logic [31:0] stage_15_out_15;
     logic [31:0] stage_15_out_16;
     logic [31:0] stage_15_out_17;
     logic [31:0] stage_15_out_18;
     logic [31:0] stage_15_out_19;
     logic [31:0] stage_15_out_20;
     logic [31:0] stage_15_out_21;
     logic [31:0] stage_15_out_22;
     logic [31:0] stage_15_out_23;
     logic [31:0] stage_15_out_24;
     logic [31:0] stage_15_out_25;
     logic [31:0] stage_15_out_26;
     logic [31:0] stage_15_out_27;
     logic [31:0] stage_15_out_28;
     logic [31:0] stage_15_out_29;
     logic [31:0] stage_15_out_30;
     logic [31:0] stage_15_out_31;
     logic [31:0] stage_15_out_32;
     logic [31:0] stage_15_out_33;
     logic [31:0] stage_15_out_34;
     logic [31:0] stage_15_out_35;
     logic [31:0] stage_15_out_36;
     logic [31:0] stage_15_out_37;
     logic [31:0] stage_15_out_38;
     logic [31:0] stage_15_out_39;
     logic [31:0] stage_15_out_40;
     logic [31:0] stage_15_out_41;
     logic [31:0] stage_15_out_42;
     logic [31:0] stage_15_out_43;
     logic [31:0] stage_15_out_44;
     logic [31:0] stage_15_out_45;
     logic [31:0] stage_15_out_46;
     logic [31:0] stage_15_out_47;
     logic [31:0] stage_15_out_48;
     logic [31:0] stage_15_out_49;
     logic [31:0] stage_15_out_50;
     logic [31:0] stage_15_out_51;
     logic [31:0] stage_15_out_52;
     logic [31:0] stage_15_out_53;
     logic [31:0] stage_15_out_54;
     logic [31:0] stage_15_out_55;
     logic [31:0] stage_15_out_56;
     logic [31:0] stage_16_out_0;
     logic [31:0] stage_16_out_1;
     logic [31:0] stage_16_out_2;
     logic [31:0] stage_16_out_3;
     logic [31:0] stage_16_out_4;
     logic [31:0] stage_16_out_5;
     logic [31:0] stage_16_out_6;
     logic [31:0] stage_16_out_7;
     logic [31:0] stage_16_out_8;
     logic [31:0] stage_16_out_9;
     logic [31:0] stage_16_out_10;
     logic [31:0] stage_16_out_11;
     logic [31:0] stage_16_out_12;
     logic [31:0] stage_16_out_13;
     logic [31:0] stage_16_out_14;
     logic [31:0] stage_16_out_15;
     logic [31:0] stage_16_out_16;
     logic [31:0] stage_16_out_17;
     logic [31:0] stage_16_out_18;
     logic [31:0] stage_16_out_19;
     logic [31:0] stage_16_out_20;
     logic [31:0] stage_16_out_21;
     logic [31:0] stage_16_out_22;
     logic [31:0] stage_16_out_23;
     logic [31:0] stage_16_out_24;
     logic [31:0] stage_16_out_25;
     logic [31:0] stage_16_out_26;
     logic [31:0] stage_16_out_27;
     logic [31:0] stage_16_out_28;
     logic [31:0] stage_16_out_29;
     logic [31:0] stage_16_out_30;
     logic [31:0] stage_16_out_31;
     logic [31:0] stage_16_out_32;
     logic [31:0] stage_16_out_33;
     logic [31:0] stage_16_out_34;
     logic [31:0] stage_16_out_35;
     logic [31:0] stage_16_out_36;
     logic [31:0] stage_16_out_37;
     logic [31:0] stage_16_out_38;
     logic [31:0] stage_16_out_39;
     logic [31:0] stage_16_out_40;
     logic [31:0] stage_16_out_41;
     logic [31:0] stage_16_out_42;
     logic [31:0] stage_16_out_43;
     logic [31:0] stage_16_out_44;
     logic [31:0] stage_16_out_45;
     logic [31:0] stage_16_out_46;
     logic [31:0] stage_16_out_47;
     logic [31:0] stage_16_out_48;
     logic [31:0] stage_16_out_49;
     logic [31:0] stage_16_out_50;
     logic [31:0] stage_16_out_51;
     logic [31:0] stage_16_out_52;
     logic [31:0] stage_16_out_53;
     logic [31:0] stage_16_out_54;
     logic [31:0] stage_16_out_55;
     logic [31:0] stage_16_out_56;
     logic [31:0] stage_17_out_0;
     logic [31:0] stage_17_out_1;
     logic [31:0] stage_17_out_2;
     logic [31:0] stage_17_out_3;
     logic [31:0] stage_17_out_4;
     logic [31:0] stage_17_out_5;
     logic [31:0] stage_17_out_6;
     logic [31:0] stage_17_out_7;
     logic [31:0] stage_17_out_8;
     logic [31:0] stage_17_out_9;
     logic [31:0] stage_17_out_10;
     logic [31:0] stage_17_out_11;
     logic [31:0] stage_17_out_12;
     logic [31:0] stage_17_out_13;
     logic [31:0] stage_17_out_14;
     logic [31:0] stage_17_out_15;
     logic [31:0] stage_17_out_16;
     logic [31:0] stage_17_out_17;
     logic [31:0] stage_17_out_18;
     logic [31:0] stage_17_out_19;
     logic [31:0] stage_17_out_20;
     logic [31:0] stage_17_out_21;
     logic [31:0] stage_17_out_22;
     logic [31:0] stage_17_out_23;
     logic [31:0] stage_17_out_24;
     logic [31:0] stage_17_out_25;
     logic [31:0] stage_17_out_26;
     logic [31:0] stage_17_out_27;
     logic [31:0] stage_17_out_28;
     logic [31:0] stage_17_out_29;
     logic [31:0] stage_17_out_30;
     logic [31:0] stage_17_out_31;
     logic [31:0] stage_17_out_32;
     logic [31:0] stage_17_out_33;
     logic [31:0] stage_17_out_34;
     logic [31:0] stage_17_out_35;
     logic [31:0] stage_17_out_36;
     logic [31:0] stage_17_out_37;
     logic [31:0] stage_17_out_38;
     logic [31:0] stage_17_out_39;
     logic [31:0] stage_17_out_40;
     logic [31:0] stage_17_out_41;
     logic [31:0] stage_17_out_42;
     logic [31:0] stage_17_out_43;
     logic [31:0] stage_17_out_44;
     logic [31:0] stage_17_out_45;
     logic [31:0] stage_17_out_46;
     logic [31:0] stage_17_out_47;
     logic [31:0] stage_17_out_48;
     logic [31:0] stage_17_out_49;
     logic [31:0] stage_17_out_50;
     logic [31:0] stage_17_out_51;
     logic [31:0] stage_17_out_52;
     logic [31:0] stage_17_out_53;
     logic [31:0] stage_17_out_54;
     logic [31:0] stage_17_out_55;
     logic [31:0] stage_17_out_56;
     logic [31:0] stage_18_out_0;
     logic [31:0] stage_18_out_1;
     logic [31:0] stage_18_out_2;
     logic [31:0] stage_18_out_3;
     logic [31:0] stage_18_out_4;
     logic [31:0] stage_18_out_5;
     logic [31:0] stage_18_out_6;
     logic [31:0] stage_18_out_7;
     logic [31:0] stage_18_out_8;
     logic [31:0] stage_18_out_9;
     logic [31:0] stage_18_out_10;
     logic [31:0] stage_18_out_11;
     logic [31:0] stage_18_out_12;
     logic [31:0] stage_18_out_13;
     logic [31:0] stage_18_out_14;
     logic [31:0] stage_18_out_15;
     logic [31:0] stage_18_out_16;
     logic [31:0] stage_18_out_17;
     logic [31:0] stage_18_out_18;
     logic [31:0] stage_18_out_19;
     logic [31:0] stage_18_out_20;
     logic [31:0] stage_18_out_21;
     logic [31:0] stage_18_out_22;
     logic [31:0] stage_18_out_23;
     logic [31:0] stage_18_out_24;
     logic [31:0] stage_18_out_25;
     logic [31:0] stage_18_out_26;
     logic [31:0] stage_18_out_27;
     logic [31:0] stage_18_out_28;
     logic [31:0] stage_18_out_29;
     logic [31:0] stage_18_out_30;
     logic [31:0] stage_18_out_31;
     logic [31:0] stage_18_out_32;
     logic [31:0] stage_18_out_33;
     logic [31:0] stage_18_out_34;
     logic [31:0] stage_18_out_35;
     logic [31:0] stage_18_out_36;
     logic [31:0] stage_18_out_37;
     logic [31:0] stage_18_out_38;
     logic [31:0] stage_18_out_39;
     logic [31:0] stage_18_out_40;
     logic [31:0] stage_18_out_41;
     logic [31:0] stage_18_out_42;
     logic [31:0] stage_18_out_43;
     logic [31:0] stage_18_out_44;
     logic [31:0] stage_18_out_45;
     logic [31:0] stage_18_out_46;
     logic [31:0] stage_18_out_47;
     logic [31:0] stage_18_out_48;
     logic [31:0] stage_18_out_49;
     logic [31:0] stage_18_out_50;
     logic [31:0] stage_18_out_51;
     logic [31:0] stage_18_out_52;
     logic [31:0] stage_18_out_53;
     logic [31:0] stage_18_out_54;
     logic [31:0] stage_18_out_55;
     logic [31:0] stage_18_out_56;
     logic [31:0] stage_19_out_0;
     logic [31:0] stage_19_out_1;
     logic [31:0] stage_19_out_2;
     logic [31:0] stage_19_out_3;
     logic [31:0] stage_19_out_4;
     logic [31:0] stage_19_out_5;
     logic [31:0] stage_19_out_6;
     logic [31:0] stage_19_out_7;
     logic [31:0] stage_19_out_8;
     logic [31:0] stage_19_out_9;
     logic [31:0] stage_19_out_10;
     logic [31:0] stage_19_out_11;
     logic [31:0] stage_19_out_12;
     logic [31:0] stage_19_out_13;
     logic [31:0] stage_19_out_14;
     logic [31:0] stage_19_out_15;
     logic [31:0] stage_19_out_16;
     logic [31:0] stage_19_out_17;
     logic [31:0] stage_19_out_18;
     logic [31:0] stage_19_out_19;
     logic [31:0] stage_19_out_20;
     logic [31:0] stage_19_out_21;
     logic [31:0] stage_19_out_22;
     logic [31:0] stage_19_out_23;
     logic [31:0] stage_19_out_24;
     logic [31:0] stage_19_out_25;
     logic [31:0] stage_19_out_26;
     logic [31:0] stage_19_out_27;
     logic [31:0] stage_19_out_28;
     logic [31:0] stage_19_out_29;
     logic [31:0] stage_19_out_30;
     logic [31:0] stage_19_out_31;
     logic [31:0] stage_19_out_32;
     logic [31:0] stage_19_out_33;
     logic [31:0] stage_19_out_34;
     logic [31:0] stage_19_out_35;
     logic [31:0] stage_19_out_36;
     logic [31:0] stage_19_out_37;
     logic [31:0] stage_19_out_38;
     logic [31:0] stage_19_out_39;
     logic [31:0] stage_19_out_40;
     logic [31:0] stage_19_out_41;
     logic [31:0] stage_19_out_42;
     logic [31:0] stage_19_out_43;
     logic [31:0] stage_19_out_44;
     logic [31:0] stage_19_out_45;
     logic [31:0] stage_19_out_46;
     logic [31:0] stage_19_out_47;
     logic [31:0] stage_19_out_48;
     logic [31:0] stage_19_out_49;
     logic [31:0] stage_19_out_50;
     logic [31:0] stage_19_out_51;
     logic [31:0] stage_19_out_52;
     logic [31:0] stage_19_out_53;
     logic [31:0] stage_19_out_54;
     logic [31:0] stage_19_out_55;
     logic [31:0] stage_19_out_56;
     logic [31:0] stage_20_out_0;
     logic [31:0] stage_20_out_1;
     logic [31:0] stage_20_out_2;
     logic [31:0] stage_20_out_3;
     logic [31:0] stage_20_out_4;
     logic [31:0] stage_20_out_5;
     logic [31:0] stage_20_out_6;
     logic [31:0] stage_20_out_7;
     logic [31:0] stage_20_out_8;
     logic [31:0] stage_20_out_9;
     logic [31:0] stage_20_out_10;
     logic [31:0] stage_20_out_11;
     logic [31:0] stage_20_out_12;
     logic [31:0] stage_20_out_13;
     logic [31:0] stage_20_out_14;
     logic [31:0] stage_20_out_15;
     logic [31:0] stage_20_out_16;
     logic [31:0] stage_20_out_17;
     logic [31:0] stage_20_out_18;
     logic [31:0] stage_20_out_19;
     logic [31:0] stage_20_out_20;
     logic [31:0] stage_20_out_21;
     logic [31:0] stage_20_out_22;
     logic [31:0] stage_20_out_23;
     logic [31:0] stage_20_out_24;
     logic [31:0] stage_20_out_25;
     logic [31:0] stage_20_out_26;
     logic [31:0] stage_20_out_27;
     logic [31:0] stage_20_out_28;
     logic [31:0] stage_20_out_29;
     logic [31:0] stage_20_out_30;
     logic [31:0] stage_20_out_31;
     logic [31:0] stage_20_out_32;
     logic [31:0] stage_20_out_33;
     logic [31:0] stage_20_out_34;
     logic [31:0] stage_20_out_35;
     logic [31:0] stage_20_out_36;
     logic [31:0] stage_20_out_37;
     logic [31:0] stage_20_out_38;
     logic [31:0] stage_20_out_39;
     logic [31:0] stage_20_out_40;
     logic [31:0] stage_20_out_41;
     logic [31:0] stage_20_out_42;
     logic [31:0] stage_20_out_43;
     logic [31:0] stage_20_out_44;
     logic [31:0] stage_20_out_45;
     logic [31:0] stage_20_out_46;
     logic [31:0] stage_20_out_47;
     logic [31:0] stage_20_out_48;
     logic [31:0] stage_20_out_49;
     logic [31:0] stage_20_out_50;
     logic [31:0] stage_20_out_51;
     logic [31:0] stage_20_out_52;
     logic [31:0] stage_20_out_53;
     logic [31:0] stage_20_out_54;
     logic [31:0] stage_20_out_55;
     logic [31:0] stage_20_out_56;
     logic [31:0] stage_21_out_0;
     logic [31:0] stage_21_out_1;
     logic [31:0] stage_21_out_2;
     logic [31:0] stage_21_out_3;
     logic [31:0] stage_21_out_4;
     logic [31:0] stage_21_out_5;
     logic [31:0] stage_21_out_6;
     logic [31:0] stage_21_out_7;
     logic [31:0] stage_21_out_8;
     logic [31:0] stage_21_out_9;
     logic [31:0] stage_21_out_10;
     logic [31:0] stage_21_out_11;
     logic [31:0] stage_21_out_12;
     logic [31:0] stage_21_out_13;
     logic [31:0] stage_21_out_14;
     logic [31:0] stage_21_out_15;
     logic [31:0] stage_21_out_16;
     logic [31:0] stage_21_out_17;
     logic [31:0] stage_21_out_18;
     logic [31:0] stage_21_out_19;
     logic [31:0] stage_21_out_20;
     logic [31:0] stage_21_out_21;
     logic [31:0] stage_21_out_22;
     logic [31:0] stage_21_out_23;
     logic [31:0] stage_21_out_24;
     logic [31:0] stage_21_out_25;
     logic [31:0] stage_21_out_26;
     logic [31:0] stage_21_out_27;
     logic [31:0] stage_21_out_28;
     logic [31:0] stage_21_out_29;
     logic [31:0] stage_21_out_30;
     logic [31:0] stage_21_out_31;
     logic [31:0] stage_21_out_32;
     logic [31:0] stage_21_out_33;
     logic [31:0] stage_21_out_34;
     logic [31:0] stage_21_out_35;
     logic [31:0] stage_21_out_36;
     logic [31:0] stage_21_out_37;
     logic [31:0] stage_21_out_38;
     logic [31:0] stage_21_out_39;
     logic [31:0] stage_21_out_40;
     logic [31:0] stage_21_out_41;
     logic [31:0] stage_21_out_42;
     logic [31:0] stage_21_out_43;
     logic [31:0] stage_21_out_44;
     logic [31:0] stage_21_out_45;
     logic [31:0] stage_21_out_46;
     logic [31:0] stage_21_out_47;
     logic [31:0] stage_21_out_48;
     logic [31:0] stage_21_out_49;
     logic [31:0] stage_21_out_50;
     logic [31:0] stage_21_out_51;
     logic [31:0] stage_21_out_52;
     logic [31:0] stage_21_out_53;
     logic [31:0] stage_21_out_54;
     logic [31:0] stage_21_out_55;
     logic [31:0] stage_21_out_56;
     logic [31:0] stage_22_out_0;
     logic [31:0] stage_22_out_1;
     logic [31:0] stage_22_out_2;
     logic [31:0] stage_22_out_3;
     logic [31:0] stage_22_out_4;
     logic [31:0] stage_22_out_5;
     logic [31:0] stage_22_out_6;
     logic [31:0] stage_22_out_7;
     logic [31:0] stage_22_out_8;
     logic [31:0] stage_22_out_9;
     logic [31:0] stage_22_out_10;
     logic [31:0] stage_22_out_11;
     logic [31:0] stage_22_out_12;
     logic [31:0] stage_22_out_13;
     logic [31:0] stage_22_out_14;
     logic [31:0] stage_22_out_15;
     logic [31:0] stage_22_out_16;
     logic [31:0] stage_22_out_17;
     logic [31:0] stage_22_out_18;
     logic [31:0] stage_22_out_19;
     logic [31:0] stage_22_out_20;
     logic [31:0] stage_22_out_21;
     logic [31:0] stage_22_out_22;
     logic [31:0] stage_22_out_23;
     logic [31:0] stage_22_out_24;
     logic [31:0] stage_22_out_25;
     logic [31:0] stage_22_out_26;
     logic [31:0] stage_22_out_27;
     logic [31:0] stage_22_out_28;
     logic [31:0] stage_22_out_29;
     logic [31:0] stage_22_out_30;
     logic [31:0] stage_22_out_31;
     logic [31:0] stage_22_out_32;
     logic [31:0] stage_22_out_33;
     logic [31:0] stage_22_out_34;
     logic [31:0] stage_22_out_35;
     logic [31:0] stage_22_out_36;
     logic [31:0] stage_22_out_37;
     logic [31:0] stage_22_out_38;
     logic [31:0] stage_22_out_39;
     logic [31:0] stage_22_out_40;
     logic [31:0] stage_22_out_41;
     logic [31:0] stage_22_out_42;
     logic [31:0] stage_22_out_43;
     logic [31:0] stage_22_out_44;
     logic [31:0] stage_22_out_45;
     logic [31:0] stage_22_out_46;
     logic [31:0] stage_22_out_47;
     logic [31:0] stage_22_out_48;
     logic [31:0] stage_22_out_49;
     logic [31:0] stage_22_out_50;
     logic [31:0] stage_22_out_51;
     logic [31:0] stage_22_out_52;
     logic [31:0] stage_22_out_53;
     logic [31:0] stage_22_out_54;
     logic [31:0] stage_22_out_55;
     logic [31:0] stage_22_out_56;
     logic [31:0] stage_23_out_0;
     logic [31:0] stage_23_out_1;
     logic [31:0] stage_23_out_2;
     logic [31:0] stage_23_out_3;
     logic [31:0] stage_23_out_4;
     logic [31:0] stage_23_out_5;
     logic [31:0] stage_23_out_6;
     logic [31:0] stage_23_out_7;
     logic [31:0] stage_23_out_8;
     logic [31:0] stage_23_out_9;
     logic [31:0] stage_23_out_10;
     logic [31:0] stage_23_out_11;
     logic [31:0] stage_23_out_12;
     logic [31:0] stage_23_out_13;
     logic [31:0] stage_23_out_14;
     logic [31:0] stage_23_out_15;
     logic [31:0] stage_23_out_16;
     logic [31:0] stage_23_out_17;
     logic [31:0] stage_23_out_18;
     logic [31:0] stage_23_out_19;
     logic [31:0] stage_23_out_20;
     logic [31:0] stage_23_out_21;
     logic [31:0] stage_23_out_22;
     logic [31:0] stage_23_out_23;
     logic [31:0] stage_23_out_24;
     logic [31:0] stage_23_out_25;
     logic [31:0] stage_23_out_26;
     logic [31:0] stage_23_out_27;
     logic [31:0] stage_23_out_28;
     logic [31:0] stage_23_out_29;
     logic [31:0] stage_23_out_30;
     logic [31:0] stage_23_out_31;
     logic [31:0] stage_23_out_32;
     logic [31:0] stage_23_out_33;
     logic [31:0] stage_23_out_34;
     logic [31:0] stage_23_out_35;
     logic [31:0] stage_23_out_36;
     logic [31:0] stage_23_out_37;
     logic [31:0] stage_23_out_38;
     logic [31:0] stage_23_out_39;
     logic [31:0] stage_23_out_40;
     logic [31:0] stage_23_out_41;
     logic [31:0] stage_23_out_42;
     logic [31:0] stage_23_out_43;
     logic [31:0] stage_23_out_44;
     logic [31:0] stage_23_out_45;
     logic [31:0] stage_23_out_46;
     logic [31:0] stage_23_out_47;
     logic [31:0] stage_23_out_48;
     logic [31:0] stage_23_out_49;
     logic [31:0] stage_23_out_50;
     logic [31:0] stage_23_out_51;
     logic [31:0] stage_23_out_52;
     logic [31:0] stage_23_out_53;
     logic [31:0] stage_23_out_54;
     logic [31:0] stage_23_out_55;
     logic [31:0] stage_23_out_56;
     logic [31:0] stage_24_out_0;
     logic [31:0] stage_24_out_1;
     logic [31:0] stage_24_out_2;
     logic [31:0] stage_24_out_3;
     logic [31:0] stage_24_out_4;
     logic [31:0] stage_24_out_5;
     logic [31:0] stage_24_out_6;
     logic [31:0] stage_24_out_7;
     logic [31:0] stage_24_out_8;
     logic [31:0] stage_24_out_9;
     logic [31:0] stage_24_out_10;
     logic [31:0] stage_24_out_11;
     logic [31:0] stage_24_out_12;
     logic [31:0] stage_24_out_13;
     logic [31:0] stage_24_out_14;
     logic [31:0] stage_24_out_15;
     logic [31:0] stage_24_out_16;
     logic [31:0] stage_24_out_17;
     logic [31:0] stage_24_out_18;
     logic [31:0] stage_24_out_19;
     logic [31:0] stage_24_out_20;
     logic [31:0] stage_24_out_21;
     logic [31:0] stage_24_out_22;
     logic [31:0] stage_24_out_23;
     logic [31:0] stage_24_out_24;
     logic [31:0] stage_24_out_25;
     logic [31:0] stage_24_out_26;
     logic [31:0] stage_24_out_27;
     logic [31:0] stage_24_out_28;
     logic [31:0] stage_24_out_29;
     logic [31:0] stage_24_out_30;
     logic [31:0] stage_24_out_31;
     logic [31:0] stage_24_out_32;
     logic [31:0] stage_24_out_33;
     logic [31:0] stage_24_out_34;
     logic [31:0] stage_24_out_35;
     logic [31:0] stage_24_out_36;
     logic [31:0] stage_24_out_37;
     logic [31:0] stage_24_out_38;
     logic [31:0] stage_24_out_39;
     logic [31:0] stage_24_out_40;
     logic [31:0] stage_24_out_41;
     logic [31:0] stage_24_out_42;
     logic [31:0] stage_24_out_43;
     logic [31:0] stage_24_out_44;
     logic [31:0] stage_24_out_45;
     logic [31:0] stage_24_out_46;
     logic [31:0] stage_24_out_47;
     logic [31:0] stage_24_out_48;
     logic [31:0] stage_24_out_49;
     logic [31:0] stage_24_out_50;
     logic [31:0] stage_24_out_51;
     logic [31:0] stage_24_out_52;
     logic [31:0] stage_24_out_53;
     logic [31:0] stage_24_out_54;
     logic [31:0] stage_24_out_55;
     logic [31:0] stage_24_out_56;
     logic [31:0] stage_25_out_0;
     logic [31:0] stage_25_out_1;
     logic [31:0] stage_25_out_2;
     logic [31:0] stage_25_out_3;
     logic [31:0] stage_25_out_4;
     logic [31:0] stage_25_out_5;
     logic [31:0] stage_25_out_6;
     logic [31:0] stage_25_out_7;
     logic [31:0] stage_25_out_8;
     logic [31:0] stage_25_out_9;
     logic [31:0] stage_25_out_10;
     logic [31:0] stage_25_out_11;
     logic [31:0] stage_25_out_12;
     logic [31:0] stage_25_out_13;
     logic [31:0] stage_25_out_14;
     logic [31:0] stage_25_out_15;
     logic [31:0] stage_25_out_16;
     logic [31:0] stage_25_out_17;
     logic [31:0] stage_25_out_18;
     logic [31:0] stage_25_out_19;
     logic [31:0] stage_25_out_20;
     logic [31:0] stage_25_out_21;
     logic [31:0] stage_25_out_22;
     logic [31:0] stage_25_out_23;
     logic [31:0] stage_25_out_24;
     logic [31:0] stage_25_out_25;
     logic [31:0] stage_25_out_26;
     logic [31:0] stage_25_out_27;
     logic [31:0] stage_25_out_28;
     logic [31:0] stage_25_out_29;
     logic [31:0] stage_25_out_30;
     logic [31:0] stage_25_out_31;
     logic [31:0] stage_25_out_32;
     logic [31:0] stage_25_out_33;
     logic [31:0] stage_25_out_34;
     logic [31:0] stage_25_out_35;
     logic [31:0] stage_25_out_36;
     logic [31:0] stage_25_out_37;
     logic [31:0] stage_25_out_38;
     logic [31:0] stage_25_out_39;
     logic [31:0] stage_25_out_40;
     logic [31:0] stage_25_out_41;
     logic [31:0] stage_25_out_42;
     logic [31:0] stage_25_out_43;
     logic [31:0] stage_25_out_44;
     logic [31:0] stage_25_out_45;
     logic [31:0] stage_25_out_46;
     logic [31:0] stage_25_out_47;
     logic [31:0] stage_25_out_48;
     logic [31:0] stage_25_out_49;
     logic [31:0] stage_25_out_50;
     logic [31:0] stage_25_out_51;
     logic [31:0] stage_25_out_52;
     logic [31:0] stage_25_out_53;
     logic [31:0] stage_25_out_54;
     logic [31:0] stage_25_out_55;
     logic [31:0] stage_25_out_56;
    assign stage_0_out_1 = (data_1 <= data_2) ? data_1 : data_2;
    assign stage_0_out_2 = (data_1 <= data_2) ? data_2 : data_1;
    assign stage_0_out_4 = (data_4 <= data_6) ? data_4 : data_6;
    assign stage_0_out_6 = (data_4 <= data_6) ? data_6 : data_4;
    assign stage_0_out_5 = (data_5 <= data_7) ? data_5 : data_7;
    assign stage_0_out_7 = (data_5 <= data_7) ? data_7 : data_5;
    assign stage_0_out_8 = (data_8 <= data_10) ? data_8 : data_10;
    assign stage_0_out_10 = (data_8 <= data_10) ? data_10 : data_8;
    assign stage_0_out_9 = (data_9 <= data_11) ? data_9 : data_11;
    assign stage_0_out_11 = (data_9 <= data_11) ? data_11 : data_9;
    assign stage_0_out_12 = (data_12 <= data_14) ? data_12 : data_14;
    assign stage_0_out_14 = (data_12 <= data_14) ? data_14 : data_12;
    assign stage_0_out_13 = (data_13 <= data_15) ? data_13 : data_15;
    assign stage_0_out_15 = (data_13 <= data_15) ? data_15 : data_13;
    assign stage_0_out_16 = (data_16 <= data_18) ? data_16 : data_18;
    assign stage_0_out_18 = (data_16 <= data_18) ? data_18 : data_16;
    assign stage_0_out_17 = (data_17 <= data_19) ? data_17 : data_19;
    assign stage_0_out_19 = (data_17 <= data_19) ? data_19 : data_17;
    assign stage_0_out_20 = (data_20 <= data_22) ? data_20 : data_22;
    assign stage_0_out_22 = (data_20 <= data_22) ? data_22 : data_20;
    assign stage_0_out_21 = (data_21 <= data_23) ? data_21 : data_23;
    assign stage_0_out_23 = (data_21 <= data_23) ? data_23 : data_21;
    assign stage_0_out_24 = (data_24 <= data_26) ? data_24 : data_26;
    assign stage_0_out_26 = (data_24 <= data_26) ? data_26 : data_24;
    assign stage_0_out_25 = (data_25 <= data_27) ? data_25 : data_27;
    assign stage_0_out_27 = (data_25 <= data_27) ? data_27 : data_25;
    assign stage_0_out_28 = (data_28 <= data_30) ? data_28 : data_30;
    assign stage_0_out_30 = (data_28 <= data_30) ? data_30 : data_28;
    assign stage_0_out_29 = (data_29 <= data_31) ? data_29 : data_31;
    assign stage_0_out_31 = (data_29 <= data_31) ? data_31 : data_29;
    assign stage_0_out_32 = (data_32 <= data_34) ? data_32 : data_34;
    assign stage_0_out_34 = (data_32 <= data_34) ? data_34 : data_32;
    assign stage_0_out_33 = (data_33 <= data_35) ? data_33 : data_35;
    assign stage_0_out_35 = (data_33 <= data_35) ? data_35 : data_33;
    assign stage_0_out_36 = (data_36 <= data_38) ? data_36 : data_38;
    assign stage_0_out_38 = (data_36 <= data_38) ? data_38 : data_36;
    assign stage_0_out_37 = (data_37 <= data_39) ? data_37 : data_39;
    assign stage_0_out_39 = (data_37 <= data_39) ? data_39 : data_37;
    assign stage_0_out_40 = (data_40 <= data_42) ? data_40 : data_42;
    assign stage_0_out_42 = (data_40 <= data_42) ? data_42 : data_40;
    assign stage_0_out_41 = (data_41 <= data_43) ? data_41 : data_43;
    assign stage_0_out_43 = (data_41 <= data_43) ? data_43 : data_41;
    assign stage_0_out_44 = (data_44 <= data_46) ? data_44 : data_46;
    assign stage_0_out_46 = (data_44 <= data_46) ? data_46 : data_44;
    assign stage_0_out_45 = (data_45 <= data_47) ? data_45 : data_47;
    assign stage_0_out_47 = (data_45 <= data_47) ? data_47 : data_45;
    assign stage_0_out_48 = (data_48 <= data_50) ? data_48 : data_50;
    assign stage_0_out_50 = (data_48 <= data_50) ? data_50 : data_48;
    assign stage_0_out_49 = (data_49 <= data_51) ? data_49 : data_51;
    assign stage_0_out_51 = (data_49 <= data_51) ? data_51 : data_49;
    assign stage_0_out_52 = (data_52 <= data_54) ? data_52 : data_54;
    assign stage_0_out_54 = (data_52 <= data_54) ? data_54 : data_52;
    assign stage_0_out_0 = (data_0 <= data_3) ? data_0 : data_3;
    assign stage_0_out_3 = (data_0 <= data_3) ? data_3 : data_0;
    assign stage_0_out_53 = data_53;
    assign stage_0_out_55 = data_55;
    assign stage_0_out_56 = data_56;
    assign stage_1_out_2 = (stage_0_out_2 <= stage_0_out_3) ? stage_0_out_2 : stage_0_out_3;
    assign stage_1_out_3 = (stage_0_out_2 <= stage_0_out_3) ? stage_0_out_3 : stage_0_out_2;
    assign stage_1_out_4 = (stage_0_out_4 <= stage_0_out_5) ? stage_0_out_4 : stage_0_out_5;
    assign stage_1_out_5 = (stage_0_out_4 <= stage_0_out_5) ? stage_0_out_5 : stage_0_out_4;
    assign stage_1_out_6 = (stage_0_out_6 <= stage_0_out_7) ? stage_0_out_6 : stage_0_out_7;
    assign stage_1_out_7 = (stage_0_out_6 <= stage_0_out_7) ? stage_0_out_7 : stage_0_out_6;
    assign stage_1_out_8 = (stage_0_out_8 <= stage_0_out_9) ? stage_0_out_8 : stage_0_out_9;
    assign stage_1_out_9 = (stage_0_out_8 <= stage_0_out_9) ? stage_0_out_9 : stage_0_out_8;
    assign stage_1_out_10 = (stage_0_out_10 <= stage_0_out_11) ? stage_0_out_10 : stage_0_out_11;
    assign stage_1_out_11 = (stage_0_out_10 <= stage_0_out_11) ? stage_0_out_11 : stage_0_out_10;
    assign stage_1_out_12 = (stage_0_out_12 <= stage_0_out_13) ? stage_0_out_12 : stage_0_out_13;
    assign stage_1_out_13 = (stage_0_out_12 <= stage_0_out_13) ? stage_0_out_13 : stage_0_out_12;
    assign stage_1_out_14 = (stage_0_out_14 <= stage_0_out_15) ? stage_0_out_14 : stage_0_out_15;
    assign stage_1_out_15 = (stage_0_out_14 <= stage_0_out_15) ? stage_0_out_15 : stage_0_out_14;
    assign stage_1_out_16 = (stage_0_out_16 <= stage_0_out_17) ? stage_0_out_16 : stage_0_out_17;
    assign stage_1_out_17 = (stage_0_out_16 <= stage_0_out_17) ? stage_0_out_17 : stage_0_out_16;
    assign stage_1_out_18 = (stage_0_out_18 <= stage_0_out_19) ? stage_0_out_18 : stage_0_out_19;
    assign stage_1_out_19 = (stage_0_out_18 <= stage_0_out_19) ? stage_0_out_19 : stage_0_out_18;
    assign stage_1_out_20 = (stage_0_out_20 <= stage_0_out_21) ? stage_0_out_20 : stage_0_out_21;
    assign stage_1_out_21 = (stage_0_out_20 <= stage_0_out_21) ? stage_0_out_21 : stage_0_out_20;
    assign stage_1_out_22 = (stage_0_out_22 <= stage_0_out_23) ? stage_0_out_22 : stage_0_out_23;
    assign stage_1_out_23 = (stage_0_out_22 <= stage_0_out_23) ? stage_0_out_23 : stage_0_out_22;
    assign stage_1_out_24 = (stage_0_out_24 <= stage_0_out_25) ? stage_0_out_24 : stage_0_out_25;
    assign stage_1_out_25 = (stage_0_out_24 <= stage_0_out_25) ? stage_0_out_25 : stage_0_out_24;
    assign stage_1_out_26 = (stage_0_out_26 <= stage_0_out_27) ? stage_0_out_26 : stage_0_out_27;
    assign stage_1_out_27 = (stage_0_out_26 <= stage_0_out_27) ? stage_0_out_27 : stage_0_out_26;
    assign stage_1_out_28 = (stage_0_out_28 <= stage_0_out_29) ? stage_0_out_28 : stage_0_out_29;
    assign stage_1_out_29 = (stage_0_out_28 <= stage_0_out_29) ? stage_0_out_29 : stage_0_out_28;
    assign stage_1_out_30 = (stage_0_out_30 <= stage_0_out_31) ? stage_0_out_30 : stage_0_out_31;
    assign stage_1_out_31 = (stage_0_out_30 <= stage_0_out_31) ? stage_0_out_31 : stage_0_out_30;
    assign stage_1_out_32 = (stage_0_out_32 <= stage_0_out_33) ? stage_0_out_32 : stage_0_out_33;
    assign stage_1_out_33 = (stage_0_out_32 <= stage_0_out_33) ? stage_0_out_33 : stage_0_out_32;
    assign stage_1_out_34 = (stage_0_out_34 <= stage_0_out_35) ? stage_0_out_34 : stage_0_out_35;
    assign stage_1_out_35 = (stage_0_out_34 <= stage_0_out_35) ? stage_0_out_35 : stage_0_out_34;
    assign stage_1_out_36 = (stage_0_out_36 <= stage_0_out_37) ? stage_0_out_36 : stage_0_out_37;
    assign stage_1_out_37 = (stage_0_out_36 <= stage_0_out_37) ? stage_0_out_37 : stage_0_out_36;
    assign stage_1_out_38 = (stage_0_out_38 <= stage_0_out_39) ? stage_0_out_38 : stage_0_out_39;
    assign stage_1_out_39 = (stage_0_out_38 <= stage_0_out_39) ? stage_0_out_39 : stage_0_out_38;
    assign stage_1_out_40 = (stage_0_out_40 <= stage_0_out_41) ? stage_0_out_40 : stage_0_out_41;
    assign stage_1_out_41 = (stage_0_out_40 <= stage_0_out_41) ? stage_0_out_41 : stage_0_out_40;
    assign stage_1_out_42 = (stage_0_out_42 <= stage_0_out_43) ? stage_0_out_42 : stage_0_out_43;
    assign stage_1_out_43 = (stage_0_out_42 <= stage_0_out_43) ? stage_0_out_43 : stage_0_out_42;
    assign stage_1_out_44 = (stage_0_out_44 <= stage_0_out_45) ? stage_0_out_44 : stage_0_out_45;
    assign stage_1_out_45 = (stage_0_out_44 <= stage_0_out_45) ? stage_0_out_45 : stage_0_out_44;
    assign stage_1_out_46 = (stage_0_out_46 <= stage_0_out_47) ? stage_0_out_46 : stage_0_out_47;
    assign stage_1_out_47 = (stage_0_out_46 <= stage_0_out_47) ? stage_0_out_47 : stage_0_out_46;
    assign stage_1_out_48 = (stage_0_out_48 <= stage_0_out_49) ? stage_0_out_48 : stage_0_out_49;
    assign stage_1_out_49 = (stage_0_out_48 <= stage_0_out_49) ? stage_0_out_49 : stage_0_out_48;
    assign stage_1_out_50 = (stage_0_out_50 <= stage_0_out_51) ? stage_0_out_50 : stage_0_out_51;
    assign stage_1_out_51 = (stage_0_out_50 <= stage_0_out_51) ? stage_0_out_51 : stage_0_out_50;
    assign stage_1_out_52 = (stage_0_out_52 <= stage_0_out_53) ? stage_0_out_52 : stage_0_out_53;
    assign stage_1_out_53 = (stage_0_out_52 <= stage_0_out_53) ? stage_0_out_53 : stage_0_out_52;
    assign stage_1_out_0 = stage_0_out_0;
    assign stage_1_out_1 = stage_0_out_1;
    assign stage_1_out_54 = stage_0_out_54;
    assign stage_1_out_55 = stage_0_out_55;
    assign stage_1_out_56 = stage_0_out_56;
    assign stage_2_out_0 = (stage_1_out_0 <= stage_1_out_7) ? stage_1_out_0 : stage_1_out_7;
    assign stage_2_out_7 = (stage_1_out_0 <= stage_1_out_7) ? stage_1_out_7 : stage_1_out_0;
    assign stage_2_out_3 = (stage_1_out_3 <= stage_1_out_11) ? stage_1_out_3 : stage_1_out_11;
    assign stage_2_out_11 = (stage_1_out_3 <= stage_1_out_11) ? stage_1_out_11 : stage_1_out_3;
    assign stage_2_out_4 = (stage_1_out_4 <= stage_1_out_8) ? stage_1_out_4 : stage_1_out_8;
    assign stage_2_out_8 = (stage_1_out_4 <= stage_1_out_8) ? stage_1_out_8 : stage_1_out_4;
    assign stage_2_out_5 = (stage_1_out_5 <= stage_1_out_6) ? stage_1_out_5 : stage_1_out_6;
    assign stage_2_out_6 = (stage_1_out_5 <= stage_1_out_6) ? stage_1_out_6 : stage_1_out_5;
    assign stage_2_out_9 = (stage_1_out_9 <= stage_1_out_10) ? stage_1_out_9 : stage_1_out_10;
    assign stage_2_out_10 = (stage_1_out_9 <= stage_1_out_10) ? stage_1_out_10 : stage_1_out_9;
    assign stage_2_out_12 = (stage_1_out_12 <= stage_1_out_20) ? stage_1_out_12 : stage_1_out_20;
    assign stage_2_out_20 = (stage_1_out_12 <= stage_1_out_20) ? stage_1_out_20 : stage_1_out_12;
    assign stage_2_out_13 = (stage_1_out_13 <= stage_1_out_14) ? stage_1_out_13 : stage_1_out_14;
    assign stage_2_out_14 = (stage_1_out_13 <= stage_1_out_14) ? stage_1_out_14 : stage_1_out_13;
    assign stage_2_out_15 = (stage_1_out_15 <= stage_1_out_23) ? stage_1_out_15 : stage_1_out_23;
    assign stage_2_out_23 = (stage_1_out_15 <= stage_1_out_23) ? stage_1_out_23 : stage_1_out_15;
    assign stage_2_out_16 = (stage_1_out_16 <= stage_1_out_24) ? stage_1_out_16 : stage_1_out_24;
    assign stage_2_out_24 = (stage_1_out_16 <= stage_1_out_24) ? stage_1_out_24 : stage_1_out_16;
    assign stage_2_out_17 = (stage_1_out_17 <= stage_1_out_18) ? stage_1_out_17 : stage_1_out_18;
    assign stage_2_out_18 = (stage_1_out_17 <= stage_1_out_18) ? stage_1_out_18 : stage_1_out_17;
    assign stage_2_out_19 = (stage_1_out_19 <= stage_1_out_27) ? stage_1_out_19 : stage_1_out_27;
    assign stage_2_out_27 = (stage_1_out_19 <= stage_1_out_27) ? stage_1_out_27 : stage_1_out_19;
    assign stage_2_out_21 = (stage_1_out_21 <= stage_1_out_22) ? stage_1_out_21 : stage_1_out_22;
    assign stage_2_out_22 = (stage_1_out_21 <= stage_1_out_22) ? stage_1_out_22 : stage_1_out_21;
    assign stage_2_out_25 = (stage_1_out_25 <= stage_1_out_26) ? stage_1_out_25 : stage_1_out_26;
    assign stage_2_out_26 = (stage_1_out_25 <= stage_1_out_26) ? stage_1_out_26 : stage_1_out_25;
    assign stage_2_out_28 = (stage_1_out_28 <= stage_1_out_36) ? stage_1_out_28 : stage_1_out_36;
    assign stage_2_out_36 = (stage_1_out_28 <= stage_1_out_36) ? stage_1_out_36 : stage_1_out_28;
    assign stage_2_out_29 = (stage_1_out_29 <= stage_1_out_30) ? stage_1_out_29 : stage_1_out_30;
    assign stage_2_out_30 = (stage_1_out_29 <= stage_1_out_30) ? stage_1_out_30 : stage_1_out_29;
    assign stage_2_out_31 = (stage_1_out_31 <= stage_1_out_39) ? stage_1_out_31 : stage_1_out_39;
    assign stage_2_out_39 = (stage_1_out_31 <= stage_1_out_39) ? stage_1_out_39 : stage_1_out_31;
    assign stage_2_out_32 = (stage_1_out_32 <= stage_1_out_40) ? stage_1_out_32 : stage_1_out_40;
    assign stage_2_out_40 = (stage_1_out_32 <= stage_1_out_40) ? stage_1_out_40 : stage_1_out_32;
    assign stage_2_out_33 = (stage_1_out_33 <= stage_1_out_34) ? stage_1_out_33 : stage_1_out_34;
    assign stage_2_out_34 = (stage_1_out_33 <= stage_1_out_34) ? stage_1_out_34 : stage_1_out_33;
    assign stage_2_out_35 = (stage_1_out_35 <= stage_1_out_43) ? stage_1_out_35 : stage_1_out_43;
    assign stage_2_out_43 = (stage_1_out_35 <= stage_1_out_43) ? stage_1_out_43 : stage_1_out_35;
    assign stage_2_out_37 = (stage_1_out_37 <= stage_1_out_38) ? stage_1_out_37 : stage_1_out_38;
    assign stage_2_out_38 = (stage_1_out_37 <= stage_1_out_38) ? stage_1_out_38 : stage_1_out_37;
    assign stage_2_out_41 = (stage_1_out_41 <= stage_1_out_42) ? stage_1_out_41 : stage_1_out_42;
    assign stage_2_out_42 = (stage_1_out_41 <= stage_1_out_42) ? stage_1_out_42 : stage_1_out_41;
    assign stage_2_out_44 = (stage_1_out_44 <= stage_1_out_52) ? stage_1_out_44 : stage_1_out_52;
    assign stage_2_out_52 = (stage_1_out_44 <= stage_1_out_52) ? stage_1_out_52 : stage_1_out_44;
    assign stage_2_out_45 = (stage_1_out_45 <= stage_1_out_46) ? stage_1_out_45 : stage_1_out_46;
    assign stage_2_out_46 = (stage_1_out_45 <= stage_1_out_46) ? stage_1_out_46 : stage_1_out_45;
    assign stage_2_out_47 = (stage_1_out_47 <= stage_1_out_51) ? stage_1_out_47 : stage_1_out_51;
    assign stage_2_out_51 = (stage_1_out_47 <= stage_1_out_51) ? stage_1_out_51 : stage_1_out_47;
    assign stage_2_out_48 = (stage_1_out_48 <= stage_1_out_55) ? stage_1_out_48 : stage_1_out_55;
    assign stage_2_out_55 = (stage_1_out_48 <= stage_1_out_55) ? stage_1_out_55 : stage_1_out_48;
    assign stage_2_out_49 = (stage_1_out_49 <= stage_1_out_50) ? stage_1_out_49 : stage_1_out_50;
    assign stage_2_out_50 = (stage_1_out_49 <= stage_1_out_50) ? stage_1_out_50 : stage_1_out_49;
    assign stage_2_out_53 = (stage_1_out_53 <= stage_1_out_54) ? stage_1_out_53 : stage_1_out_54;
    assign stage_2_out_54 = (stage_1_out_53 <= stage_1_out_54) ? stage_1_out_54 : stage_1_out_53;
    assign stage_2_out_1 = stage_1_out_1;
    assign stage_2_out_2 = stage_1_out_2;
    assign stage_2_out_56 = stage_1_out_56;
    assign stage_3_out_1 = (stage_2_out_1 <= stage_2_out_9) ? stage_2_out_1 : stage_2_out_9;
    assign stage_3_out_9 = (stage_2_out_1 <= stage_2_out_9) ? stage_2_out_9 : stage_2_out_1;
    assign stage_3_out_2 = (stage_2_out_2 <= stage_2_out_10) ? stage_2_out_2 : stage_2_out_10;
    assign stage_3_out_10 = (stage_2_out_2 <= stage_2_out_10) ? stage_2_out_10 : stage_2_out_2;
    assign stage_3_out_7 = (stage_2_out_7 <= stage_2_out_11) ? stage_2_out_7 : stage_2_out_11;
    assign stage_3_out_11 = (stage_2_out_7 <= stage_2_out_11) ? stage_2_out_11 : stage_2_out_7;
    assign stage_3_out_12 = (stage_2_out_12 <= stage_2_out_16) ? stage_2_out_12 : stage_2_out_16;
    assign stage_3_out_16 = (stage_2_out_12 <= stage_2_out_16) ? stage_2_out_16 : stage_2_out_12;
    assign stage_3_out_13 = (stage_2_out_13 <= stage_2_out_21) ? stage_2_out_13 : stage_2_out_21;
    assign stage_3_out_21 = (stage_2_out_13 <= stage_2_out_21) ? stage_2_out_21 : stage_2_out_13;
    assign stage_3_out_14 = (stage_2_out_14 <= stage_2_out_22) ? stage_2_out_14 : stage_2_out_22;
    assign stage_3_out_22 = (stage_2_out_14 <= stage_2_out_22) ? stage_2_out_22 : stage_2_out_14;
    assign stage_3_out_15 = (stage_2_out_15 <= stage_2_out_19) ? stage_2_out_15 : stage_2_out_19;
    assign stage_3_out_19 = (stage_2_out_15 <= stage_2_out_19) ? stage_2_out_19 : stage_2_out_15;
    assign stage_3_out_17 = (stage_2_out_17 <= stage_2_out_25) ? stage_2_out_17 : stage_2_out_25;
    assign stage_3_out_25 = (stage_2_out_17 <= stage_2_out_25) ? stage_2_out_25 : stage_2_out_17;
    assign stage_3_out_18 = (stage_2_out_18 <= stage_2_out_26) ? stage_2_out_18 : stage_2_out_26;
    assign stage_3_out_26 = (stage_2_out_18 <= stage_2_out_26) ? stage_2_out_26 : stage_2_out_18;
    assign stage_3_out_20 = (stage_2_out_20 <= stage_2_out_24) ? stage_2_out_20 : stage_2_out_24;
    assign stage_3_out_24 = (stage_2_out_20 <= stage_2_out_24) ? stage_2_out_24 : stage_2_out_20;
    assign stage_3_out_23 = (stage_2_out_23 <= stage_2_out_27) ? stage_2_out_23 : stage_2_out_27;
    assign stage_3_out_27 = (stage_2_out_23 <= stage_2_out_27) ? stage_2_out_27 : stage_2_out_23;
    assign stage_3_out_28 = (stage_2_out_28 <= stage_2_out_32) ? stage_2_out_28 : stage_2_out_32;
    assign stage_3_out_32 = (stage_2_out_28 <= stage_2_out_32) ? stage_2_out_32 : stage_2_out_28;
    assign stage_3_out_29 = (stage_2_out_29 <= stage_2_out_37) ? stage_2_out_29 : stage_2_out_37;
    assign stage_3_out_37 = (stage_2_out_29 <= stage_2_out_37) ? stage_2_out_37 : stage_2_out_29;
    assign stage_3_out_30 = (stage_2_out_30 <= stage_2_out_38) ? stage_2_out_30 : stage_2_out_38;
    assign stage_3_out_38 = (stage_2_out_30 <= stage_2_out_38) ? stage_2_out_38 : stage_2_out_30;
    assign stage_3_out_31 = (stage_2_out_31 <= stage_2_out_35) ? stage_2_out_31 : stage_2_out_35;
    assign stage_3_out_35 = (stage_2_out_31 <= stage_2_out_35) ? stage_2_out_35 : stage_2_out_31;
    assign stage_3_out_33 = (stage_2_out_33 <= stage_2_out_41) ? stage_2_out_33 : stage_2_out_41;
    assign stage_3_out_41 = (stage_2_out_33 <= stage_2_out_41) ? stage_2_out_41 : stage_2_out_33;
    assign stage_3_out_34 = (stage_2_out_34 <= stage_2_out_42) ? stage_2_out_34 : stage_2_out_42;
    assign stage_3_out_42 = (stage_2_out_34 <= stage_2_out_42) ? stage_2_out_42 : stage_2_out_34;
    assign stage_3_out_36 = (stage_2_out_36 <= stage_2_out_40) ? stage_2_out_36 : stage_2_out_40;
    assign stage_3_out_40 = (stage_2_out_36 <= stage_2_out_40) ? stage_2_out_40 : stage_2_out_36;
    assign stage_3_out_39 = (stage_2_out_39 <= stage_2_out_43) ? stage_2_out_39 : stage_2_out_43;
    assign stage_3_out_43 = (stage_2_out_39 <= stage_2_out_43) ? stage_2_out_43 : stage_2_out_39;
    assign stage_3_out_44 = (stage_2_out_44 <= stage_2_out_48) ? stage_2_out_44 : stage_2_out_48;
    assign stage_3_out_48 = (stage_2_out_44 <= stage_2_out_48) ? stage_2_out_48 : stage_2_out_44;
    assign stage_3_out_45 = (stage_2_out_45 <= stage_2_out_53) ? stage_2_out_45 : stage_2_out_53;
    assign stage_3_out_53 = (stage_2_out_45 <= stage_2_out_53) ? stage_2_out_53 : stage_2_out_45;
    assign stage_3_out_46 = (stage_2_out_46 <= stage_2_out_54) ? stage_2_out_46 : stage_2_out_54;
    assign stage_3_out_54 = (stage_2_out_46 <= stage_2_out_54) ? stage_2_out_54 : stage_2_out_46;
    assign stage_3_out_52 = (stage_2_out_52 <= stage_2_out_55) ? stage_2_out_52 : stage_2_out_55;
    assign stage_3_out_55 = (stage_2_out_52 <= stage_2_out_55) ? stage_2_out_55 : stage_2_out_52;
    assign stage_3_out_0 = stage_2_out_0;
    assign stage_3_out_3 = stage_2_out_3;
    assign stage_3_out_4 = stage_2_out_4;
    assign stage_3_out_5 = stage_2_out_5;
    assign stage_3_out_6 = stage_2_out_6;
    assign stage_3_out_8 = stage_2_out_8;
    assign stage_3_out_47 = stage_2_out_47;
    assign stage_3_out_49 = stage_2_out_49;
    assign stage_3_out_50 = stage_2_out_50;
    assign stage_3_out_51 = stage_2_out_51;
    assign stage_3_out_56 = stage_2_out_56;
    assign stage_4_out_0 = (stage_3_out_0 <= stage_3_out_31) ? stage_3_out_0 : stage_3_out_31;
    assign stage_4_out_31 = (stage_3_out_0 <= stage_3_out_31) ? stage_3_out_31 : stage_3_out_0;
    assign stage_4_out_3 = (stage_3_out_3 <= stage_3_out_7) ? stage_3_out_3 : stage_3_out_7;
    assign stage_4_out_7 = (stage_3_out_3 <= stage_3_out_7) ? stage_3_out_7 : stage_3_out_3;
    assign stage_4_out_5 = (stage_3_out_5 <= stage_3_out_9) ? stage_3_out_5 : stage_3_out_9;
    assign stage_4_out_9 = (stage_3_out_5 <= stage_3_out_9) ? stage_3_out_9 : stage_3_out_5;
    assign stage_4_out_6 = (stage_3_out_6 <= stage_3_out_10) ? stage_3_out_6 : stage_3_out_10;
    assign stage_4_out_10 = (stage_3_out_6 <= stage_3_out_10) ? stage_3_out_10 : stage_3_out_6;
    assign stage_4_out_8 = (stage_3_out_8 <= stage_3_out_40) ? stage_3_out_8 : stage_3_out_40;
    assign stage_4_out_40 = (stage_3_out_8 <= stage_3_out_40) ? stage_3_out_40 : stage_3_out_8;
    assign stage_4_out_11 = (stage_3_out_11 <= stage_3_out_43) ? stage_3_out_11 : stage_3_out_43;
    assign stage_4_out_43 = (stage_3_out_11 <= stage_3_out_43) ? stage_3_out_43 : stage_3_out_11;
    assign stage_4_out_12 = (stage_3_out_12 <= stage_3_out_44) ? stage_3_out_12 : stage_3_out_44;
    assign stage_4_out_44 = (stage_3_out_12 <= stage_3_out_44) ? stage_3_out_44 : stage_3_out_12;
    assign stage_4_out_13 = (stage_3_out_13 <= stage_3_out_17) ? stage_3_out_13 : stage_3_out_17;
    assign stage_4_out_17 = (stage_3_out_13 <= stage_3_out_17) ? stage_3_out_17 : stage_3_out_13;
    assign stage_4_out_14 = (stage_3_out_14 <= stage_3_out_18) ? stage_3_out_14 : stage_3_out_18;
    assign stage_4_out_18 = (stage_3_out_14 <= stage_3_out_18) ? stage_3_out_18 : stage_3_out_14;
    assign stage_4_out_15 = (stage_3_out_15 <= stage_3_out_47) ? stage_3_out_15 : stage_3_out_47;
    assign stage_4_out_47 = (stage_3_out_15 <= stage_3_out_47) ? stage_3_out_47 : stage_3_out_15;
    assign stage_4_out_16 = (stage_3_out_16 <= stage_3_out_20) ? stage_3_out_16 : stage_3_out_20;
    assign stage_4_out_20 = (stage_3_out_16 <= stage_3_out_20) ? stage_3_out_20 : stage_3_out_16;
    assign stage_4_out_19 = (stage_3_out_19 <= stage_3_out_23) ? stage_3_out_19 : stage_3_out_23;
    assign stage_4_out_23 = (stage_3_out_19 <= stage_3_out_23) ? stage_3_out_23 : stage_3_out_19;
    assign stage_4_out_21 = (stage_3_out_21 <= stage_3_out_25) ? stage_3_out_21 : stage_3_out_25;
    assign stage_4_out_25 = (stage_3_out_21 <= stage_3_out_25) ? stage_3_out_25 : stage_3_out_21;
    assign stage_4_out_22 = (stage_3_out_22 <= stage_3_out_26) ? stage_3_out_22 : stage_3_out_26;
    assign stage_4_out_26 = (stage_3_out_22 <= stage_3_out_26) ? stage_3_out_26 : stage_3_out_22;
    assign stage_4_out_24 = (stage_3_out_24 <= stage_3_out_55) ? stage_3_out_24 : stage_3_out_55;
    assign stage_4_out_55 = (stage_3_out_24 <= stage_3_out_55) ? stage_3_out_55 : stage_3_out_24;
    assign stage_4_out_29 = (stage_3_out_29 <= stage_3_out_33) ? stage_3_out_29 : stage_3_out_33;
    assign stage_4_out_33 = (stage_3_out_29 <= stage_3_out_33) ? stage_3_out_33 : stage_3_out_29;
    assign stage_4_out_30 = (stage_3_out_30 <= stage_3_out_34) ? stage_3_out_30 : stage_3_out_34;
    assign stage_4_out_34 = (stage_3_out_30 <= stage_3_out_34) ? stage_3_out_34 : stage_3_out_30;
    assign stage_4_out_32 = (stage_3_out_32 <= stage_3_out_36) ? stage_3_out_32 : stage_3_out_36;
    assign stage_4_out_36 = (stage_3_out_32 <= stage_3_out_36) ? stage_3_out_36 : stage_3_out_32;
    assign stage_4_out_35 = (stage_3_out_35 <= stage_3_out_39) ? stage_3_out_35 : stage_3_out_39;
    assign stage_4_out_39 = (stage_3_out_35 <= stage_3_out_39) ? stage_3_out_39 : stage_3_out_35;
    assign stage_4_out_37 = (stage_3_out_37 <= stage_3_out_41) ? stage_3_out_37 : stage_3_out_41;
    assign stage_4_out_41 = (stage_3_out_37 <= stage_3_out_41) ? stage_3_out_41 : stage_3_out_37;
    assign stage_4_out_38 = (stage_3_out_38 <= stage_3_out_42) ? stage_3_out_38 : stage_3_out_42;
    assign stage_4_out_42 = (stage_3_out_38 <= stage_3_out_42) ? stage_3_out_42 : stage_3_out_38;
    assign stage_4_out_45 = (stage_3_out_45 <= stage_3_out_49) ? stage_3_out_45 : stage_3_out_49;
    assign stage_4_out_49 = (stage_3_out_45 <= stage_3_out_49) ? stage_3_out_49 : stage_3_out_45;
    assign stage_4_out_46 = (stage_3_out_46 <= stage_3_out_50) ? stage_3_out_46 : stage_3_out_50;
    assign stage_4_out_50 = (stage_3_out_46 <= stage_3_out_50) ? stage_3_out_50 : stage_3_out_46;
    assign stage_4_out_48 = (stage_3_out_48 <= stage_3_out_52) ? stage_3_out_48 : stage_3_out_52;
    assign stage_4_out_52 = (stage_3_out_48 <= stage_3_out_52) ? stage_3_out_52 : stage_3_out_48;
    assign stage_4_out_27 = (stage_3_out_27 <= stage_3_out_28) ? stage_3_out_27 : stage_3_out_28;
    assign stage_4_out_28 = (stage_3_out_27 <= stage_3_out_28) ? stage_3_out_28 : stage_3_out_27;
    assign stage_4_out_1 = stage_3_out_1;
    assign stage_4_out_2 = stage_3_out_2;
    assign stage_4_out_4 = stage_3_out_4;
    assign stage_4_out_51 = stage_3_out_51;
    assign stage_4_out_53 = stage_3_out_53;
    assign stage_4_out_54 = stage_3_out_54;
    assign stage_4_out_56 = stage_3_out_56;
    assign stage_5_out_0 = (stage_4_out_0 <= stage_4_out_15) ? stage_4_out_0 : stage_4_out_15;
    assign stage_5_out_15 = (stage_4_out_0 <= stage_4_out_15) ? stage_4_out_15 : stage_4_out_0;
    assign stage_5_out_1 = (stage_4_out_1 <= stage_4_out_5) ? stage_4_out_1 : stage_4_out_5;
    assign stage_5_out_5 = (stage_4_out_1 <= stage_4_out_5) ? stage_4_out_5 : stage_4_out_1;
    assign stage_5_out_2 = (stage_4_out_2 <= stage_4_out_6) ? stage_4_out_2 : stage_4_out_6;
    assign stage_5_out_6 = (stage_4_out_2 <= stage_4_out_6) ? stage_4_out_6 : stage_4_out_2;
    assign stage_5_out_3 = (stage_4_out_3 <= stage_4_out_35) ? stage_4_out_3 : stage_4_out_35;
    assign stage_5_out_35 = (stage_4_out_3 <= stage_4_out_35) ? stage_4_out_35 : stage_4_out_3;
    assign stage_5_out_4 = (stage_4_out_4 <= stage_4_out_36) ? stage_4_out_4 : stage_4_out_36;
    assign stage_5_out_36 = (stage_4_out_4 <= stage_4_out_36) ? stage_4_out_36 : stage_4_out_4;
    assign stage_5_out_7 = (stage_4_out_7 <= stage_4_out_39) ? stage_4_out_7 : stage_4_out_39;
    assign stage_5_out_39 = (stage_4_out_7 <= stage_4_out_39) ? stage_4_out_39 : stage_4_out_7;
    assign stage_5_out_8 = (stage_4_out_8 <= stage_4_out_24) ? stage_4_out_8 : stage_4_out_24;
    assign stage_5_out_24 = (stage_4_out_8 <= stage_4_out_24) ? stage_4_out_24 : stage_4_out_8;
    assign stage_5_out_9 = (stage_4_out_9 <= stage_4_out_41) ? stage_4_out_9 : stage_4_out_41;
    assign stage_5_out_41 = (stage_4_out_9 <= stage_4_out_41) ? stage_4_out_41 : stage_4_out_9;
    assign stage_5_out_10 = (stage_4_out_10 <= stage_4_out_42) ? stage_4_out_10 : stage_4_out_42;
    assign stage_5_out_42 = (stage_4_out_10 <= stage_4_out_42) ? stage_4_out_42 : stage_4_out_10;
    assign stage_5_out_11 = (stage_4_out_11 <= stage_4_out_27) ? stage_4_out_11 : stage_4_out_27;
    assign stage_5_out_27 = (stage_4_out_11 <= stage_4_out_27) ? stage_4_out_27 : stage_4_out_11;
    assign stage_5_out_13 = (stage_4_out_13 <= stage_4_out_45) ? stage_4_out_13 : stage_4_out_45;
    assign stage_5_out_45 = (stage_4_out_13 <= stage_4_out_45) ? stage_4_out_45 : stage_4_out_13;
    assign stage_5_out_14 = (stage_4_out_14 <= stage_4_out_46) ? stage_4_out_14 : stage_4_out_46;
    assign stage_5_out_46 = (stage_4_out_14 <= stage_4_out_46) ? stage_4_out_46 : stage_4_out_14;
    assign stage_5_out_16 = (stage_4_out_16 <= stage_4_out_48) ? stage_4_out_16 : stage_4_out_48;
    assign stage_5_out_48 = (stage_4_out_16 <= stage_4_out_48) ? stage_4_out_48 : stage_4_out_16;
    assign stage_5_out_17 = (stage_4_out_17 <= stage_4_out_21) ? stage_4_out_17 : stage_4_out_21;
    assign stage_5_out_21 = (stage_4_out_17 <= stage_4_out_21) ? stage_4_out_21 : stage_4_out_17;
    assign stage_5_out_18 = (stage_4_out_18 <= stage_4_out_22) ? stage_4_out_18 : stage_4_out_22;
    assign stage_5_out_22 = (stage_4_out_18 <= stage_4_out_22) ? stage_4_out_22 : stage_4_out_18;
    assign stage_5_out_19 = (stage_4_out_19 <= stage_4_out_51) ? stage_4_out_19 : stage_4_out_51;
    assign stage_5_out_51 = (stage_4_out_19 <= stage_4_out_51) ? stage_4_out_51 : stage_4_out_19;
    assign stage_5_out_20 = (stage_4_out_20 <= stage_4_out_52) ? stage_4_out_20 : stage_4_out_52;
    assign stage_5_out_52 = (stage_4_out_20 <= stage_4_out_52) ? stage_4_out_52 : stage_4_out_20;
    assign stage_5_out_28 = (stage_4_out_28 <= stage_4_out_44) ? stage_4_out_28 : stage_4_out_44;
    assign stage_5_out_44 = (stage_4_out_28 <= stage_4_out_44) ? stage_4_out_44 : stage_4_out_28;
    assign stage_5_out_31 = (stage_4_out_31 <= stage_4_out_47) ? stage_4_out_31 : stage_4_out_47;
    assign stage_5_out_47 = (stage_4_out_31 <= stage_4_out_47) ? stage_4_out_47 : stage_4_out_31;
    assign stage_5_out_33 = (stage_4_out_33 <= stage_4_out_37) ? stage_4_out_33 : stage_4_out_37;
    assign stage_5_out_37 = (stage_4_out_33 <= stage_4_out_37) ? stage_4_out_37 : stage_4_out_33;
    assign stage_5_out_34 = (stage_4_out_34 <= stage_4_out_38) ? stage_4_out_34 : stage_4_out_38;
    assign stage_5_out_38 = (stage_4_out_34 <= stage_4_out_38) ? stage_4_out_38 : stage_4_out_34;
    assign stage_5_out_40 = (stage_4_out_40 <= stage_4_out_55) ? stage_4_out_40 : stage_4_out_55;
    assign stage_5_out_55 = (stage_4_out_40 <= stage_4_out_55) ? stage_4_out_55 : stage_4_out_40;
    assign stage_5_out_49 = (stage_4_out_49 <= stage_4_out_53) ? stage_4_out_49 : stage_4_out_53;
    assign stage_5_out_53 = (stage_4_out_49 <= stage_4_out_53) ? stage_4_out_53 : stage_4_out_49;
    assign stage_5_out_50 = (stage_4_out_50 <= stage_4_out_54) ? stage_4_out_50 : stage_4_out_54;
    assign stage_5_out_54 = (stage_4_out_50 <= stage_4_out_54) ? stage_4_out_54 : stage_4_out_50;
    assign stage_5_out_25 = (stage_4_out_25 <= stage_4_out_29) ? stage_4_out_25 : stage_4_out_29;
    assign stage_5_out_29 = (stage_4_out_25 <= stage_4_out_29) ? stage_4_out_29 : stage_4_out_25;
    assign stage_5_out_26 = (stage_4_out_26 <= stage_4_out_30) ? stage_4_out_26 : stage_4_out_30;
    assign stage_5_out_30 = (stage_4_out_26 <= stage_4_out_30) ? stage_4_out_30 : stage_4_out_26;
    assign stage_5_out_12 = stage_4_out_12;
    assign stage_5_out_23 = stage_4_out_23;
    assign stage_5_out_32 = stage_4_out_32;
    assign stage_5_out_43 = stage_4_out_43;
    assign stage_5_out_56 = stage_4_out_56;
    assign stage_6_out_1 = (stage_5_out_1 <= stage_5_out_33) ? stage_5_out_1 : stage_5_out_33;
    assign stage_6_out_33 = (stage_5_out_1 <= stage_5_out_33) ? stage_5_out_33 : stage_5_out_1;
    assign stage_6_out_2 = (stage_5_out_2 <= stage_5_out_34) ? stage_5_out_2 : stage_5_out_34;
    assign stage_6_out_34 = (stage_5_out_2 <= stage_5_out_34) ? stage_5_out_34 : stage_5_out_2;
    assign stage_6_out_3 = (stage_5_out_3 <= stage_5_out_19) ? stage_5_out_3 : stage_5_out_19;
    assign stage_6_out_19 = (stage_5_out_3 <= stage_5_out_19) ? stage_5_out_19 : stage_5_out_3;
    assign stage_6_out_4 = (stage_5_out_4 <= stage_5_out_20) ? stage_5_out_4 : stage_5_out_20;
    assign stage_6_out_20 = (stage_5_out_4 <= stage_5_out_20) ? stage_5_out_20 : stage_5_out_4;
    assign stage_6_out_5 = (stage_5_out_5 <= stage_5_out_37) ? stage_5_out_5 : stage_5_out_37;
    assign stage_6_out_37 = (stage_5_out_5 <= stage_5_out_37) ? stage_5_out_37 : stage_5_out_5;
    assign stage_6_out_6 = (stage_5_out_6 <= stage_5_out_38) ? stage_5_out_6 : stage_5_out_38;
    assign stage_6_out_38 = (stage_5_out_6 <= stage_5_out_38) ? stage_5_out_38 : stage_5_out_6;
    assign stage_6_out_7 = (stage_5_out_7 <= stage_5_out_23) ? stage_5_out_7 : stage_5_out_23;
    assign stage_6_out_23 = (stage_5_out_7 <= stage_5_out_23) ? stage_5_out_23 : stage_5_out_7;
    assign stage_6_out_9 = (stage_5_out_9 <= stage_5_out_25) ? stage_5_out_9 : stage_5_out_25;
    assign stage_6_out_25 = (stage_5_out_9 <= stage_5_out_25) ? stage_5_out_25 : stage_5_out_9;
    assign stage_6_out_10 = (stage_5_out_10 <= stage_5_out_26) ? stage_5_out_10 : stage_5_out_26;
    assign stage_6_out_26 = (stage_5_out_10 <= stage_5_out_26) ? stage_5_out_26 : stage_5_out_10;
    assign stage_6_out_12 = (stage_5_out_12 <= stage_5_out_28) ? stage_5_out_12 : stage_5_out_28;
    assign stage_6_out_28 = (stage_5_out_12 <= stage_5_out_28) ? stage_5_out_28 : stage_5_out_12;
    assign stage_6_out_15 = (stage_5_out_15 <= stage_5_out_31) ? stage_5_out_15 : stage_5_out_31;
    assign stage_6_out_31 = (stage_5_out_15 <= stage_5_out_31) ? stage_5_out_31 : stage_5_out_15;
    assign stage_6_out_17 = (stage_5_out_17 <= stage_5_out_49) ? stage_5_out_17 : stage_5_out_49;
    assign stage_6_out_49 = (stage_5_out_17 <= stage_5_out_49) ? stage_5_out_49 : stage_5_out_17;
    assign stage_6_out_18 = (stage_5_out_18 <= stage_5_out_50) ? stage_5_out_18 : stage_5_out_50;
    assign stage_6_out_50 = (stage_5_out_18 <= stage_5_out_50) ? stage_5_out_50 : stage_5_out_18;
    assign stage_6_out_21 = (stage_5_out_21 <= stage_5_out_53) ? stage_5_out_21 : stage_5_out_53;
    assign stage_6_out_53 = (stage_5_out_21 <= stage_5_out_53) ? stage_5_out_53 : stage_5_out_21;
    assign stage_6_out_22 = (stage_5_out_22 <= stage_5_out_54) ? stage_5_out_22 : stage_5_out_54;
    assign stage_6_out_54 = (stage_5_out_22 <= stage_5_out_54) ? stage_5_out_54 : stage_5_out_22;
    assign stage_6_out_24 = (stage_5_out_24 <= stage_5_out_40) ? stage_5_out_24 : stage_5_out_40;
    assign stage_6_out_40 = (stage_5_out_24 <= stage_5_out_40) ? stage_5_out_40 : stage_5_out_24;
    assign stage_6_out_27 = (stage_5_out_27 <= stage_5_out_43) ? stage_5_out_27 : stage_5_out_43;
    assign stage_6_out_43 = (stage_5_out_27 <= stage_5_out_43) ? stage_5_out_43 : stage_5_out_27;
    assign stage_6_out_29 = (stage_5_out_29 <= stage_5_out_45) ? stage_5_out_29 : stage_5_out_45;
    assign stage_6_out_45 = (stage_5_out_29 <= stage_5_out_45) ? stage_5_out_45 : stage_5_out_29;
    assign stage_6_out_30 = (stage_5_out_30 <= stage_5_out_46) ? stage_5_out_30 : stage_5_out_46;
    assign stage_6_out_46 = (stage_5_out_30 <= stage_5_out_46) ? stage_5_out_46 : stage_5_out_30;
    assign stage_6_out_32 = (stage_5_out_32 <= stage_5_out_48) ? stage_5_out_32 : stage_5_out_48;
    assign stage_6_out_48 = (stage_5_out_32 <= stage_5_out_48) ? stage_5_out_48 : stage_5_out_32;
    assign stage_6_out_35 = (stage_5_out_35 <= stage_5_out_51) ? stage_5_out_35 : stage_5_out_51;
    assign stage_6_out_51 = (stage_5_out_35 <= stage_5_out_51) ? stage_5_out_51 : stage_5_out_35;
    assign stage_6_out_36 = (stage_5_out_36 <= stage_5_out_52) ? stage_5_out_36 : stage_5_out_52;
    assign stage_6_out_52 = (stage_5_out_36 <= stage_5_out_52) ? stage_5_out_52 : stage_5_out_36;
    assign stage_6_out_11 = (stage_5_out_11 <= stage_5_out_44) ? stage_5_out_11 : stage_5_out_44;
    assign stage_6_out_44 = (stage_5_out_11 <= stage_5_out_44) ? stage_5_out_44 : stage_5_out_11;
    assign stage_6_out_0 = stage_5_out_0;
    assign stage_6_out_8 = stage_5_out_8;
    assign stage_6_out_13 = stage_5_out_13;
    assign stage_6_out_14 = stage_5_out_14;
    assign stage_6_out_16 = stage_5_out_16;
    assign stage_6_out_39 = stage_5_out_39;
    assign stage_6_out_41 = stage_5_out_41;
    assign stage_6_out_42 = stage_5_out_42;
    assign stage_6_out_47 = stage_5_out_47;
    assign stage_6_out_55 = stage_5_out_55;
    assign stage_6_out_56 = stage_5_out_56;
    assign stage_7_out_1 = (stage_6_out_1 <= stage_6_out_17) ? stage_6_out_1 : stage_6_out_17;
    assign stage_7_out_17 = (stage_6_out_1 <= stage_6_out_17) ? stage_6_out_17 : stage_6_out_1;
    assign stage_7_out_2 = (stage_6_out_2 <= stage_6_out_18) ? stage_6_out_2 : stage_6_out_18;
    assign stage_7_out_18 = (stage_6_out_2 <= stage_6_out_18) ? stage_6_out_18 : stage_6_out_2;
    assign stage_7_out_4 = (stage_6_out_4 <= stage_6_out_30) ? stage_6_out_4 : stage_6_out_30;
    assign stage_7_out_30 = (stage_6_out_4 <= stage_6_out_30) ? stage_6_out_30 : stage_6_out_4;
    assign stage_7_out_5 = (stage_6_out_5 <= stage_6_out_21) ? stage_6_out_5 : stage_6_out_21;
    assign stage_7_out_21 = (stage_6_out_5 <= stage_6_out_21) ? stage_6_out_21 : stage_6_out_5;
    assign stage_7_out_6 = (stage_6_out_6 <= stage_6_out_22) ? stage_6_out_6 : stage_6_out_22;
    assign stage_7_out_22 = (stage_6_out_6 <= stage_6_out_22) ? stage_6_out_22 : stage_6_out_6;
    assign stage_7_out_8 = (stage_6_out_8 <= stage_6_out_29) ? stage_6_out_8 : stage_6_out_29;
    assign stage_7_out_29 = (stage_6_out_8 <= stage_6_out_29) ? stage_6_out_29 : stage_6_out_8;
    assign stage_7_out_16 = (stage_6_out_16 <= stage_6_out_32) ? stage_6_out_16 : stage_6_out_32;
    assign stage_7_out_32 = (stage_6_out_16 <= stage_6_out_32) ? stage_6_out_32 : stage_6_out_16;
    assign stage_7_out_19 = (stage_6_out_19 <= stage_6_out_35) ? stage_6_out_19 : stage_6_out_35;
    assign stage_7_out_35 = (stage_6_out_19 <= stage_6_out_35) ? stage_6_out_35 : stage_6_out_19;
    assign stage_7_out_20 = (stage_6_out_20 <= stage_6_out_36) ? stage_6_out_20 : stage_6_out_36;
    assign stage_7_out_36 = (stage_6_out_20 <= stage_6_out_36) ? stage_6_out_36 : stage_6_out_20;
    assign stage_7_out_23 = (stage_6_out_23 <= stage_6_out_39) ? stage_6_out_23 : stage_6_out_39;
    assign stage_7_out_39 = (stage_6_out_23 <= stage_6_out_39) ? stage_6_out_39 : stage_6_out_23;
    assign stage_7_out_25 = (stage_6_out_25 <= stage_6_out_51) ? stage_6_out_25 : stage_6_out_51;
    assign stage_7_out_51 = (stage_6_out_25 <= stage_6_out_51) ? stage_6_out_51 : stage_6_out_25;
    assign stage_7_out_26 = (stage_6_out_26 <= stage_6_out_47) ? stage_6_out_26 : stage_6_out_47;
    assign stage_7_out_47 = (stage_6_out_26 <= stage_6_out_47) ? stage_6_out_47 : stage_6_out_26;
    assign stage_7_out_33 = (stage_6_out_33 <= stage_6_out_49) ? stage_6_out_33 : stage_6_out_49;
    assign stage_7_out_49 = (stage_6_out_33 <= stage_6_out_49) ? stage_6_out_49 : stage_6_out_33;
    assign stage_7_out_34 = (stage_6_out_34 <= stage_6_out_50) ? stage_6_out_34 : stage_6_out_50;
    assign stage_7_out_50 = (stage_6_out_34 <= stage_6_out_50) ? stage_6_out_50 : stage_6_out_34;
    assign stage_7_out_37 = (stage_6_out_37 <= stage_6_out_53) ? stage_6_out_37 : stage_6_out_53;
    assign stage_7_out_53 = (stage_6_out_37 <= stage_6_out_53) ? stage_6_out_53 : stage_6_out_37;
    assign stage_7_out_38 = (stage_6_out_38 <= stage_6_out_54) ? stage_6_out_38 : stage_6_out_54;
    assign stage_7_out_54 = (stage_6_out_38 <= stage_6_out_54) ? stage_6_out_54 : stage_6_out_38;
    assign stage_7_out_7 = (stage_6_out_7 <= stage_6_out_44) ? stage_6_out_7 : stage_6_out_44;
    assign stage_7_out_44 = (stage_6_out_7 <= stage_6_out_44) ? stage_6_out_44 : stage_6_out_7;
    assign stage_7_out_11 = (stage_6_out_11 <= stage_6_out_48) ? stage_6_out_11 : stage_6_out_48;
    assign stage_7_out_48 = (stage_6_out_11 <= stage_6_out_48) ? stage_6_out_48 : stage_6_out_11;
    assign stage_7_out_10 = (stage_6_out_10 <= stage_6_out_27) ? stage_6_out_10 : stage_6_out_27;
    assign stage_7_out_27 = (stage_6_out_10 <= stage_6_out_27) ? stage_6_out_27 : stage_6_out_10;
    assign stage_7_out_28 = (stage_6_out_28 <= stage_6_out_45) ? stage_6_out_28 : stage_6_out_45;
    assign stage_7_out_45 = (stage_6_out_28 <= stage_6_out_45) ? stage_6_out_45 : stage_6_out_28;
    assign stage_7_out_0 = stage_6_out_0;
    assign stage_7_out_3 = stage_6_out_3;
    assign stage_7_out_9 = stage_6_out_9;
    assign stage_7_out_12 = stage_6_out_12;
    assign stage_7_out_13 = stage_6_out_13;
    assign stage_7_out_14 = stage_6_out_14;
    assign stage_7_out_15 = stage_6_out_15;
    assign stage_7_out_24 = stage_6_out_24;
    assign stage_7_out_31 = stage_6_out_31;
    assign stage_7_out_40 = stage_6_out_40;
    assign stage_7_out_41 = stage_6_out_41;
    assign stage_7_out_42 = stage_6_out_42;
    assign stage_7_out_43 = stage_6_out_43;
    assign stage_7_out_46 = stage_6_out_46;
    assign stage_7_out_52 = stage_6_out_52;
    assign stage_7_out_55 = stage_6_out_55;
    assign stage_7_out_56 = stage_6_out_56;
    assign stage_8_out_0 = (stage_7_out_0 <= stage_7_out_20) ? stage_7_out_0 : stage_7_out_20;
    assign stage_8_out_20 = (stage_7_out_0 <= stage_7_out_20) ? stage_7_out_20 : stage_7_out_0;
    assign stage_8_out_2 = (stage_7_out_2 <= stage_7_out_44) ? stage_7_out_2 : stage_7_out_44;
    assign stage_8_out_44 = (stage_7_out_2 <= stage_7_out_44) ? stage_7_out_44 : stage_7_out_2;
    assign stage_8_out_5 = (stage_7_out_5 <= stage_7_out_32) ? stage_7_out_5 : stage_7_out_32;
    assign stage_8_out_32 = (stage_7_out_5 <= stage_7_out_32) ? stage_7_out_32 : stage_7_out_5;
    assign stage_8_out_6 = (stage_7_out_6 <= stage_7_out_15) ? stage_7_out_6 : stage_7_out_15;
    assign stage_8_out_15 = (stage_7_out_6 <= stage_7_out_15) ? stage_7_out_15 : stage_7_out_6;
    assign stage_8_out_10 = (stage_7_out_10 <= stage_7_out_19) ? stage_7_out_10 : stage_7_out_19;
    assign stage_8_out_19 = (stage_7_out_10 <= stage_7_out_19) ? stage_7_out_19 : stage_7_out_10;
    assign stage_8_out_11 = (stage_7_out_11 <= stage_7_out_53) ? stage_7_out_11 : stage_7_out_53;
    assign stage_8_out_53 = (stage_7_out_11 <= stage_7_out_53) ? stage_7_out_53 : stage_7_out_11;
    assign stage_8_out_14 = (stage_7_out_14 <= stage_7_out_30) ? stage_7_out_14 : stage_7_out_30;
    assign stage_8_out_30 = (stage_7_out_14 <= stage_7_out_30) ? stage_7_out_30 : stage_7_out_14;
    assign stage_8_out_17 = (stage_7_out_17 <= stage_7_out_33) ? stage_7_out_17 : stage_7_out_33;
    assign stage_8_out_33 = (stage_7_out_17 <= stage_7_out_33) ? stage_7_out_33 : stage_7_out_17;
    assign stage_8_out_18 = (stage_7_out_18 <= stage_7_out_34) ? stage_7_out_18 : stage_7_out_34;
    assign stage_8_out_34 = (stage_7_out_18 <= stage_7_out_34) ? stage_7_out_34 : stage_7_out_18;
    assign stage_8_out_21 = (stage_7_out_21 <= stage_7_out_37) ? stage_7_out_21 : stage_7_out_37;
    assign stage_8_out_37 = (stage_7_out_21 <= stage_7_out_37) ? stage_7_out_37 : stage_7_out_21;
    assign stage_8_out_22 = (stage_7_out_22 <= stage_7_out_38) ? stage_7_out_22 : stage_7_out_38;
    assign stage_8_out_38 = (stage_7_out_22 <= stage_7_out_38) ? stage_7_out_38 : stage_7_out_22;
    assign stage_8_out_23 = (stage_7_out_23 <= stage_7_out_50) ? stage_7_out_23 : stage_7_out_50;
    assign stage_8_out_50 = (stage_7_out_23 <= stage_7_out_50) ? stage_7_out_50 : stage_7_out_23;
    assign stage_8_out_25 = (stage_7_out_25 <= stage_7_out_41) ? stage_7_out_25 : stage_7_out_41;
    assign stage_8_out_41 = (stage_7_out_25 <= stage_7_out_41) ? stage_7_out_41 : stage_7_out_25;
    assign stage_8_out_35 = (stage_7_out_35 <= stage_7_out_55) ? stage_7_out_35 : stage_7_out_55;
    assign stage_8_out_55 = (stage_7_out_35 <= stage_7_out_55) ? stage_7_out_55 : stage_7_out_35;
    assign stage_8_out_36 = (stage_7_out_36 <= stage_7_out_45) ? stage_7_out_36 : stage_7_out_45;
    assign stage_8_out_45 = (stage_7_out_36 <= stage_7_out_45) ? stage_7_out_45 : stage_7_out_36;
    assign stage_8_out_40 = (stage_7_out_40 <= stage_7_out_49) ? stage_7_out_40 : stage_7_out_49;
    assign stage_8_out_49 = (stage_7_out_40 <= stage_7_out_49) ? stage_7_out_49 : stage_7_out_40;
    assign stage_8_out_13 = (stage_7_out_13 <= stage_7_out_29) ? stage_7_out_13 : stage_7_out_29;
    assign stage_8_out_29 = (stage_7_out_13 <= stage_7_out_29) ? stage_7_out_29 : stage_7_out_13;
    assign stage_8_out_26 = (stage_7_out_26 <= stage_7_out_42) ? stage_7_out_26 : stage_7_out_42;
    assign stage_8_out_42 = (stage_7_out_26 <= stage_7_out_42) ? stage_7_out_42 : stage_7_out_26;
    assign stage_8_out_28 = (stage_7_out_28 <= stage_7_out_56) ? stage_7_out_28 : stage_7_out_56;
    assign stage_8_out_56 = (stage_7_out_28 <= stage_7_out_56) ? stage_7_out_56 : stage_7_out_28;
    assign stage_8_out_1 = stage_7_out_1;
    assign stage_8_out_3 = stage_7_out_3;
    assign stage_8_out_4 = stage_7_out_4;
    assign stage_8_out_7 = stage_7_out_7;
    assign stage_8_out_8 = stage_7_out_8;
    assign stage_8_out_9 = stage_7_out_9;
    assign stage_8_out_12 = stage_7_out_12;
    assign stage_8_out_16 = stage_7_out_16;
    assign stage_8_out_24 = stage_7_out_24;
    assign stage_8_out_27 = stage_7_out_27;
    assign stage_8_out_31 = stage_7_out_31;
    assign stage_8_out_39 = stage_7_out_39;
    assign stage_8_out_43 = stage_7_out_43;
    assign stage_8_out_46 = stage_7_out_46;
    assign stage_8_out_47 = stage_7_out_47;
    assign stage_8_out_48 = stage_7_out_48;
    assign stage_8_out_51 = stage_7_out_51;
    assign stage_8_out_52 = stage_7_out_52;
    assign stage_8_out_54 = stage_7_out_54;
    assign stage_9_out_3 = (stage_8_out_3 <= stage_8_out_21) ? stage_8_out_3 : stage_8_out_21;
    assign stage_9_out_21 = (stage_8_out_3 <= stage_8_out_21) ? stage_8_out_21 : stage_8_out_3;
    assign stage_9_out_7 = (stage_8_out_7 <= stage_8_out_25) ? stage_8_out_7 : stage_8_out_25;
    assign stage_9_out_25 = (stage_8_out_7 <= stage_8_out_25) ? stage_8_out_25 : stage_8_out_7;
    assign stage_9_out_9 = (stage_8_out_9 <= stage_8_out_18) ? stage_8_out_9 : stage_8_out_18;
    assign stage_9_out_18 = (stage_8_out_9 <= stage_8_out_18) ? stage_8_out_18 : stage_8_out_9;
    assign stage_9_out_11 = (stage_8_out_11 <= stage_8_out_35) ? stage_8_out_11 : stage_8_out_35;
    assign stage_9_out_35 = (stage_8_out_11 <= stage_8_out_35) ? stage_8_out_35 : stage_8_out_11;
    assign stage_9_out_14 = (stage_8_out_14 <= stage_8_out_32) ? stage_8_out_14 : stage_8_out_32;
    assign stage_9_out_32 = (stage_8_out_14 <= stage_8_out_32) ? stage_8_out_32 : stage_8_out_14;
    assign stage_9_out_20 = (stage_8_out_20 <= stage_8_out_44) ? stage_8_out_20 : stage_8_out_44;
    assign stage_9_out_44 = (stage_8_out_20 <= stage_8_out_44) ? stage_8_out_44 : stage_8_out_20;
    assign stage_9_out_22 = (stage_8_out_22 <= stage_8_out_31) ? stage_8_out_22 : stage_8_out_31;
    assign stage_9_out_31 = (stage_8_out_22 <= stage_8_out_31) ? stage_8_out_31 : stage_8_out_22;
    assign stage_9_out_23 = (stage_8_out_23 <= stage_8_out_41) ? stage_8_out_23 : stage_8_out_41;
    assign stage_9_out_41 = (stage_8_out_23 <= stage_8_out_41) ? stage_8_out_41 : stage_8_out_23;
    assign stage_9_out_24 = (stage_8_out_24 <= stage_8_out_33) ? stage_8_out_24 : stage_8_out_33;
    assign stage_9_out_33 = (stage_8_out_24 <= stage_8_out_33) ? stage_8_out_33 : stage_8_out_24;
    assign stage_9_out_30 = (stage_8_out_30 <= stage_8_out_48) ? stage_8_out_30 : stage_8_out_48;
    assign stage_9_out_48 = (stage_8_out_30 <= stage_8_out_48) ? stage_8_out_48 : stage_8_out_30;
    assign stage_9_out_34 = (stage_8_out_34 <= stage_8_out_52) ? stage_8_out_34 : stage_8_out_52;
    assign stage_9_out_52 = (stage_8_out_34 <= stage_8_out_52) ? stage_8_out_52 : stage_8_out_34;
    assign stage_9_out_37 = (stage_8_out_37 <= stage_8_out_46) ? stage_8_out_37 : stage_8_out_46;
    assign stage_9_out_46 = (stage_8_out_37 <= stage_8_out_46) ? stage_8_out_46 : stage_8_out_37;
    assign stage_9_out_15 = (stage_8_out_15 <= stage_8_out_36) ? stage_8_out_15 : stage_8_out_36;
    assign stage_9_out_36 = (stage_8_out_15 <= stage_8_out_36) ? stage_8_out_36 : stage_8_out_15;
    assign stage_9_out_19 = (stage_8_out_19 <= stage_8_out_40) ? stage_8_out_19 : stage_8_out_40;
    assign stage_9_out_40 = (stage_8_out_19 <= stage_8_out_40) ? stage_8_out_40 : stage_8_out_19;
    assign stage_9_out_17 = (stage_8_out_17 <= stage_8_out_29) ? stage_8_out_17 : stage_8_out_29;
    assign stage_9_out_29 = (stage_8_out_17 <= stage_8_out_29) ? stage_8_out_29 : stage_8_out_17;
    assign stage_9_out_26 = (stage_8_out_26 <= stage_8_out_38) ? stage_8_out_26 : stage_8_out_38;
    assign stage_9_out_38 = (stage_8_out_26 <= stage_8_out_38) ? stage_8_out_38 : stage_8_out_26;
    assign stage_9_out_0 = stage_8_out_0;
    assign stage_9_out_1 = stage_8_out_1;
    assign stage_9_out_2 = stage_8_out_2;
    assign stage_9_out_4 = stage_8_out_4;
    assign stage_9_out_5 = stage_8_out_5;
    assign stage_9_out_6 = stage_8_out_6;
    assign stage_9_out_8 = stage_8_out_8;
    assign stage_9_out_10 = stage_8_out_10;
    assign stage_9_out_12 = stage_8_out_12;
    assign stage_9_out_13 = stage_8_out_13;
    assign stage_9_out_16 = stage_8_out_16;
    assign stage_9_out_27 = stage_8_out_27;
    assign stage_9_out_28 = stage_8_out_28;
    assign stage_9_out_39 = stage_8_out_39;
    assign stage_9_out_42 = stage_8_out_42;
    assign stage_9_out_43 = stage_8_out_43;
    assign stage_9_out_45 = stage_8_out_45;
    assign stage_9_out_47 = stage_8_out_47;
    assign stage_9_out_49 = stage_8_out_49;
    assign stage_9_out_50 = stage_8_out_50;
    assign stage_9_out_51 = stage_8_out_51;
    assign stage_9_out_53 = stage_8_out_53;
    assign stage_9_out_54 = stage_8_out_54;
    assign stage_9_out_55 = stage_8_out_55;
    assign stage_9_out_56 = stage_8_out_56;
    assign stage_10_out_3 = (stage_9_out_3 <= stage_9_out_30) ? stage_9_out_3 : stage_9_out_30;
    assign stage_10_out_30 = (stage_9_out_3 <= stage_9_out_30) ? stage_9_out_30 : stage_9_out_3;
    assign stage_10_out_6 = (stage_9_out_6 <= stage_9_out_24) ? stage_9_out_6 : stage_9_out_24;
    assign stage_10_out_24 = (stage_9_out_6 <= stage_9_out_24) ? stage_9_out_24 : stage_9_out_6;
    assign stage_10_out_7 = (stage_9_out_7 <= stage_9_out_34) ? stage_9_out_7 : stage_9_out_34;
    assign stage_10_out_34 = (stage_9_out_7 <= stage_9_out_34) ? stage_9_out_34 : stage_9_out_7;
    assign stage_10_out_9 = (stage_9_out_9 <= stage_9_out_36) ? stage_9_out_9 : stage_9_out_36;
    assign stage_10_out_36 = (stage_9_out_9 <= stage_9_out_36) ? stage_9_out_36 : stage_9_out_9;
    assign stage_10_out_10 = (stage_9_out_10 <= stage_9_out_37) ? stage_9_out_10 : stage_9_out_37;
    assign stage_10_out_37 = (stage_9_out_10 <= stage_9_out_37) ? stage_9_out_37 : stage_9_out_10;
    assign stage_10_out_15 = (stage_9_out_15 <= stage_9_out_33) ? stage_9_out_15 : stage_9_out_33;
    assign stage_10_out_33 = (stage_9_out_15 <= stage_9_out_33) ? stage_9_out_33 : stage_9_out_15;
    assign stage_10_out_18 = (stage_9_out_18 <= stage_9_out_45) ? stage_9_out_18 : stage_9_out_45;
    assign stage_10_out_45 = (stage_9_out_18 <= stage_9_out_45) ? stage_9_out_45 : stage_9_out_18;
    assign stage_10_out_19 = (stage_9_out_19 <= stage_9_out_46) ? stage_9_out_19 : stage_9_out_46;
    assign stage_10_out_46 = (stage_9_out_19 <= stage_9_out_46) ? stage_9_out_46 : stage_9_out_19;
    assign stage_10_out_20 = (stage_9_out_20 <= stage_9_out_29) ? stage_9_out_20 : stage_9_out_29;
    assign stage_10_out_29 = (stage_9_out_20 <= stage_9_out_29) ? stage_9_out_29 : stage_9_out_20;
    assign stage_10_out_21 = (stage_9_out_21 <= stage_9_out_48) ? stage_9_out_21 : stage_9_out_48;
    assign stage_10_out_48 = (stage_9_out_21 <= stage_9_out_48) ? stage_9_out_48 : stage_9_out_21;
    assign stage_10_out_22 = (stage_9_out_22 <= stage_9_out_40) ? stage_9_out_22 : stage_9_out_40;
    assign stage_10_out_40 = (stage_9_out_22 <= stage_9_out_40) ? stage_9_out_40 : stage_9_out_22;
    assign stage_10_out_25 = (stage_9_out_25 <= stage_9_out_52) ? stage_9_out_25 : stage_9_out_52;
    assign stage_10_out_52 = (stage_9_out_25 <= stage_9_out_52) ? stage_9_out_52 : stage_9_out_25;
    assign stage_10_out_26 = (stage_9_out_26 <= stage_9_out_35) ? stage_9_out_26 : stage_9_out_35;
    assign stage_10_out_35 = (stage_9_out_26 <= stage_9_out_35) ? stage_9_out_35 : stage_9_out_26;
    assign stage_10_out_31 = (stage_9_out_31 <= stage_9_out_49) ? stage_9_out_31 : stage_9_out_49;
    assign stage_10_out_49 = (stage_9_out_31 <= stage_9_out_49) ? stage_9_out_49 : stage_9_out_31;
    assign stage_10_out_23 = (stage_9_out_23 <= stage_9_out_28) ? stage_9_out_23 : stage_9_out_28;
    assign stage_10_out_28 = (stage_9_out_23 <= stage_9_out_28) ? stage_9_out_28 : stage_9_out_23;
    assign stage_10_out_27 = (stage_9_out_27 <= stage_9_out_32) ? stage_9_out_27 : stage_9_out_32;
    assign stage_10_out_32 = (stage_9_out_27 <= stage_9_out_32) ? stage_9_out_32 : stage_9_out_27;
    assign stage_10_out_0 = stage_9_out_0;
    assign stage_10_out_1 = stage_9_out_1;
    assign stage_10_out_2 = stage_9_out_2;
    assign stage_10_out_4 = stage_9_out_4;
    assign stage_10_out_5 = stage_9_out_5;
    assign stage_10_out_8 = stage_9_out_8;
    assign stage_10_out_11 = stage_9_out_11;
    assign stage_10_out_12 = stage_9_out_12;
    assign stage_10_out_13 = stage_9_out_13;
    assign stage_10_out_14 = stage_9_out_14;
    assign stage_10_out_16 = stage_9_out_16;
    assign stage_10_out_17 = stage_9_out_17;
    assign stage_10_out_38 = stage_9_out_38;
    assign stage_10_out_39 = stage_9_out_39;
    assign stage_10_out_41 = stage_9_out_41;
    assign stage_10_out_42 = stage_9_out_42;
    assign stage_10_out_43 = stage_9_out_43;
    assign stage_10_out_44 = stage_9_out_44;
    assign stage_10_out_47 = stage_9_out_47;
    assign stage_10_out_50 = stage_9_out_50;
    assign stage_10_out_51 = stage_9_out_51;
    assign stage_10_out_53 = stage_9_out_53;
    assign stage_10_out_54 = stage_9_out_54;
    assign stage_10_out_55 = stage_9_out_55;
    assign stage_10_out_56 = stage_9_out_56;
    assign stage_11_out_10 = (stage_10_out_10 <= stage_10_out_22) ? stage_10_out_10 : stage_10_out_22;
    assign stage_11_out_22 = (stage_10_out_10 <= stage_10_out_22) ? stage_10_out_22 : stage_10_out_10;
    assign stage_11_out_18 = (stage_10_out_18 <= stage_10_out_24) ? stage_10_out_18 : stage_10_out_24;
    assign stage_11_out_24 = (stage_10_out_18 <= stage_10_out_24) ? stage_10_out_24 : stage_10_out_18;
    assign stage_11_out_31 = (stage_10_out_31 <= stage_10_out_37) ? stage_10_out_31 : stage_10_out_37;
    assign stage_11_out_37 = (stage_10_out_31 <= stage_10_out_37) ? stage_10_out_37 : stage_10_out_31;
    assign stage_11_out_33 = (stage_10_out_33 <= stage_10_out_45) ? stage_10_out_33 : stage_10_out_45;
    assign stage_11_out_45 = (stage_10_out_33 <= stage_10_out_45) ? stage_10_out_45 : stage_10_out_33;
    assign stage_11_out_7 = (stage_10_out_7 <= stage_10_out_32) ? stage_10_out_7 : stage_10_out_32;
    assign stage_11_out_32 = (stage_10_out_7 <= stage_10_out_32) ? stage_10_out_32 : stage_10_out_7;
    assign stage_11_out_19 = (stage_10_out_19 <= stage_10_out_34) ? stage_10_out_19 : stage_10_out_34;
    assign stage_11_out_34 = (stage_10_out_19 <= stage_10_out_34) ? stage_10_out_34 : stage_10_out_19;
    assign stage_11_out_21 = (stage_10_out_21 <= stage_10_out_36) ? stage_10_out_21 : stage_10_out_36;
    assign stage_11_out_36 = (stage_10_out_21 <= stage_10_out_36) ? stage_10_out_36 : stage_10_out_21;
    assign stage_11_out_23 = (stage_10_out_23 <= stage_10_out_48) ? stage_10_out_23 : stage_10_out_48;
    assign stage_11_out_48 = (stage_10_out_23 <= stage_10_out_48) ? stage_10_out_48 : stage_10_out_23;
    assign stage_11_out_11 = (stage_10_out_11 <= stage_10_out_26) ? stage_10_out_11 : stage_10_out_26;
    assign stage_11_out_26 = (stage_10_out_11 <= stage_10_out_26) ? stage_10_out_26 : stage_10_out_11;
    assign stage_11_out_29 = (stage_10_out_29 <= stage_10_out_44) ? stage_10_out_29 : stage_10_out_44;
    assign stage_11_out_44 = (stage_10_out_29 <= stage_10_out_44) ? stage_10_out_44 : stage_10_out_29;
    assign stage_11_out_0 = stage_10_out_0;
    assign stage_11_out_1 = stage_10_out_1;
    assign stage_11_out_2 = stage_10_out_2;
    assign stage_11_out_3 = stage_10_out_3;
    assign stage_11_out_4 = stage_10_out_4;
    assign stage_11_out_5 = stage_10_out_5;
    assign stage_11_out_6 = stage_10_out_6;
    assign stage_11_out_8 = stage_10_out_8;
    assign stage_11_out_9 = stage_10_out_9;
    assign stage_11_out_12 = stage_10_out_12;
    assign stage_11_out_13 = stage_10_out_13;
    assign stage_11_out_14 = stage_10_out_14;
    assign stage_11_out_15 = stage_10_out_15;
    assign stage_11_out_16 = stage_10_out_16;
    assign stage_11_out_17 = stage_10_out_17;
    assign stage_11_out_20 = stage_10_out_20;
    assign stage_11_out_25 = stage_10_out_25;
    assign stage_11_out_27 = stage_10_out_27;
    assign stage_11_out_28 = stage_10_out_28;
    assign stage_11_out_30 = stage_10_out_30;
    assign stage_11_out_35 = stage_10_out_35;
    assign stage_11_out_38 = stage_10_out_38;
    assign stage_11_out_39 = stage_10_out_39;
    assign stage_11_out_40 = stage_10_out_40;
    assign stage_11_out_41 = stage_10_out_41;
    assign stage_11_out_42 = stage_10_out_42;
    assign stage_11_out_43 = stage_10_out_43;
    assign stage_11_out_46 = stage_10_out_46;
    assign stage_11_out_47 = stage_10_out_47;
    assign stage_11_out_49 = stage_10_out_49;
    assign stage_11_out_50 = stage_10_out_50;
    assign stage_11_out_51 = stage_10_out_51;
    assign stage_11_out_52 = stage_10_out_52;
    assign stage_11_out_53 = stage_10_out_53;
    assign stage_11_out_54 = stage_10_out_54;
    assign stage_11_out_55 = stage_10_out_55;
    assign stage_11_out_56 = stage_10_out_56;
    assign stage_12_out_22 = (stage_11_out_22 <= stage_11_out_29) ? stage_11_out_22 : stage_11_out_29;
    assign stage_12_out_29 = (stage_11_out_22 <= stage_11_out_29) ? stage_11_out_29 : stage_11_out_22;
    assign stage_12_out_24 = (stage_11_out_24 <= stage_11_out_30) ? stage_11_out_24 : stage_11_out_30;
    assign stage_12_out_30 = (stage_11_out_24 <= stage_11_out_30) ? stage_11_out_30 : stage_11_out_24;
    assign stage_12_out_25 = (stage_11_out_25 <= stage_11_out_31) ? stage_11_out_25 : stage_11_out_31;
    assign stage_12_out_31 = (stage_11_out_25 <= stage_11_out_31) ? stage_11_out_31 : stage_11_out_25;
    assign stage_12_out_26 = (stage_11_out_26 <= stage_11_out_33) ? stage_11_out_26 : stage_11_out_33;
    assign stage_12_out_33 = (stage_11_out_26 <= stage_11_out_33) ? stage_11_out_33 : stage_11_out_26;
    assign stage_12_out_18 = (stage_11_out_18 <= stage_11_out_21) ? stage_11_out_18 : stage_11_out_21;
    assign stage_12_out_21 = (stage_11_out_18 <= stage_11_out_21) ? stage_11_out_21 : stage_11_out_18;
    assign stage_12_out_34 = (stage_11_out_34 <= stage_11_out_37) ? stage_11_out_34 : stage_11_out_37;
    assign stage_12_out_37 = (stage_11_out_34 <= stage_11_out_37) ? stage_11_out_37 : stage_11_out_34;
    assign stage_12_out_11 = (stage_11_out_11 <= stage_11_out_19) ? stage_11_out_11 : stage_11_out_19;
    assign stage_12_out_19 = (stage_11_out_11 <= stage_11_out_19) ? stage_11_out_19 : stage_11_out_11;
    assign stage_12_out_36 = (stage_11_out_36 <= stage_11_out_44) ? stage_11_out_36 : stage_11_out_44;
    assign stage_12_out_44 = (stage_11_out_36 <= stage_11_out_44) ? stage_11_out_44 : stage_11_out_36;
    assign stage_12_out_0 = stage_11_out_0;
    assign stage_12_out_1 = stage_11_out_1;
    assign stage_12_out_2 = stage_11_out_2;
    assign stage_12_out_3 = stage_11_out_3;
    assign stage_12_out_4 = stage_11_out_4;
    assign stage_12_out_5 = stage_11_out_5;
    assign stage_12_out_6 = stage_11_out_6;
    assign stage_12_out_7 = stage_11_out_7;
    assign stage_12_out_8 = stage_11_out_8;
    assign stage_12_out_9 = stage_11_out_9;
    assign stage_12_out_10 = stage_11_out_10;
    assign stage_12_out_12 = stage_11_out_12;
    assign stage_12_out_13 = stage_11_out_13;
    assign stage_12_out_14 = stage_11_out_14;
    assign stage_12_out_15 = stage_11_out_15;
    assign stage_12_out_16 = stage_11_out_16;
    assign stage_12_out_17 = stage_11_out_17;
    assign stage_12_out_20 = stage_11_out_20;
    assign stage_12_out_23 = stage_11_out_23;
    assign stage_12_out_27 = stage_11_out_27;
    assign stage_12_out_28 = stage_11_out_28;
    assign stage_12_out_32 = stage_11_out_32;
    assign stage_12_out_35 = stage_11_out_35;
    assign stage_12_out_38 = stage_11_out_38;
    assign stage_12_out_39 = stage_11_out_39;
    assign stage_12_out_40 = stage_11_out_40;
    assign stage_12_out_41 = stage_11_out_41;
    assign stage_12_out_42 = stage_11_out_42;
    assign stage_12_out_43 = stage_11_out_43;
    assign stage_12_out_45 = stage_11_out_45;
    assign stage_12_out_46 = stage_11_out_46;
    assign stage_12_out_47 = stage_11_out_47;
    assign stage_12_out_48 = stage_11_out_48;
    assign stage_12_out_49 = stage_11_out_49;
    assign stage_12_out_50 = stage_11_out_50;
    assign stage_12_out_51 = stage_11_out_51;
    assign stage_12_out_52 = stage_11_out_52;
    assign stage_12_out_53 = stage_11_out_53;
    assign stage_12_out_54 = stage_11_out_54;
    assign stage_12_out_55 = stage_11_out_55;
    assign stage_12_out_56 = stage_11_out_56;
    assign stage_13_out_19 = (stage_12_out_19 <= stage_12_out_25) ? stage_12_out_19 : stage_12_out_25;
    assign stage_13_out_25 = (stage_12_out_19 <= stage_12_out_25) ? stage_12_out_25 : stage_12_out_19;
    assign stage_13_out_22 = (stage_12_out_22 <= stage_12_out_32) ? stage_12_out_22 : stage_12_out_32;
    assign stage_13_out_32 = (stage_12_out_22 <= stage_12_out_32) ? stage_12_out_32 : stage_12_out_22;
    assign stage_13_out_23 = (stage_12_out_23 <= stage_12_out_33) ? stage_12_out_23 : stage_12_out_33;
    assign stage_13_out_33 = (stage_12_out_23 <= stage_12_out_33) ? stage_12_out_33 : stage_12_out_23;
    assign stage_13_out_30 = (stage_12_out_30 <= stage_12_out_36) ? stage_12_out_30 : stage_12_out_36;
    assign stage_13_out_36 = (stage_12_out_30 <= stage_12_out_36) ? stage_12_out_36 : stage_12_out_30;
    assign stage_13_out_15 = (stage_12_out_15 <= stage_12_out_21) ? stage_12_out_15 : stage_12_out_21;
    assign stage_13_out_21 = (stage_12_out_15 <= stage_12_out_21) ? stage_12_out_21 : stage_12_out_15;
    assign stage_13_out_34 = (stage_12_out_34 <= stage_12_out_40) ? stage_12_out_34 : stage_12_out_40;
    assign stage_13_out_40 = (stage_12_out_34 <= stage_12_out_40) ? stage_12_out_40 : stage_12_out_34;
    assign stage_13_out_26 = (stage_12_out_26 <= stage_12_out_28) ? stage_12_out_26 : stage_12_out_28;
    assign stage_13_out_28 = (stage_12_out_26 <= stage_12_out_28) ? stage_12_out_28 : stage_12_out_26;
    assign stage_13_out_27 = (stage_12_out_27 <= stage_12_out_29) ? stage_12_out_27 : stage_12_out_29;
    assign stage_13_out_29 = (stage_12_out_27 <= stage_12_out_29) ? stage_12_out_29 : stage_12_out_27;
    assign stage_13_out_0 = stage_12_out_0;
    assign stage_13_out_1 = stage_12_out_1;
    assign stage_13_out_2 = stage_12_out_2;
    assign stage_13_out_3 = stage_12_out_3;
    assign stage_13_out_4 = stage_12_out_4;
    assign stage_13_out_5 = stage_12_out_5;
    assign stage_13_out_6 = stage_12_out_6;
    assign stage_13_out_7 = stage_12_out_7;
    assign stage_13_out_8 = stage_12_out_8;
    assign stage_13_out_9 = stage_12_out_9;
    assign stage_13_out_10 = stage_12_out_10;
    assign stage_13_out_11 = stage_12_out_11;
    assign stage_13_out_12 = stage_12_out_12;
    assign stage_13_out_13 = stage_12_out_13;
    assign stage_13_out_14 = stage_12_out_14;
    assign stage_13_out_16 = stage_12_out_16;
    assign stage_13_out_17 = stage_12_out_17;
    assign stage_13_out_18 = stage_12_out_18;
    assign stage_13_out_20 = stage_12_out_20;
    assign stage_13_out_24 = stage_12_out_24;
    assign stage_13_out_31 = stage_12_out_31;
    assign stage_13_out_35 = stage_12_out_35;
    assign stage_13_out_37 = stage_12_out_37;
    assign stage_13_out_38 = stage_12_out_38;
    assign stage_13_out_39 = stage_12_out_39;
    assign stage_13_out_41 = stage_12_out_41;
    assign stage_13_out_42 = stage_12_out_42;
    assign stage_13_out_43 = stage_12_out_43;
    assign stage_13_out_44 = stage_12_out_44;
    assign stage_13_out_45 = stage_12_out_45;
    assign stage_13_out_46 = stage_12_out_46;
    assign stage_13_out_47 = stage_12_out_47;
    assign stage_13_out_48 = stage_12_out_48;
    assign stage_13_out_49 = stage_12_out_49;
    assign stage_13_out_50 = stage_12_out_50;
    assign stage_13_out_51 = stage_12_out_51;
    assign stage_13_out_52 = stage_12_out_52;
    assign stage_13_out_53 = stage_12_out_53;
    assign stage_13_out_54 = stage_12_out_54;
    assign stage_13_out_55 = stage_12_out_55;
    assign stage_13_out_56 = stage_12_out_56;
    assign stage_14_out_21 = (stage_13_out_21 <= stage_13_out_24) ? stage_13_out_21 : stage_13_out_24;
    assign stage_14_out_24 = (stage_13_out_21 <= stage_13_out_24) ? stage_13_out_24 : stage_13_out_21;
    assign stage_14_out_31 = (stage_13_out_31 <= stage_13_out_34) ? stage_13_out_31 : stage_13_out_34;
    assign stage_14_out_34 = (stage_13_out_31 <= stage_13_out_34) ? stage_13_out_34 : stage_13_out_31;
    assign stage_14_out_11 = (stage_13_out_11 <= stage_13_out_29) ? stage_13_out_11 : stage_13_out_29;
    assign stage_14_out_29 = (stage_13_out_11 <= stage_13_out_29) ? stage_13_out_29 : stage_13_out_11;
    assign stage_14_out_26 = (stage_13_out_26 <= stage_13_out_44) ? stage_13_out_26 : stage_13_out_44;
    assign stage_14_out_44 = (stage_13_out_26 <= stage_13_out_44) ? stage_13_out_44 : stage_13_out_26;
    assign stage_14_out_19 = (stage_13_out_19 <= stage_13_out_30) ? stage_13_out_19 : stage_13_out_30;
    assign stage_14_out_30 = (stage_13_out_19 <= stage_13_out_30) ? stage_13_out_30 : stage_13_out_19;
    assign stage_14_out_25 = (stage_13_out_25 <= stage_13_out_36) ? stage_13_out_25 : stage_13_out_36;
    assign stage_14_out_36 = (stage_13_out_25 <= stage_13_out_36) ? stage_13_out_36 : stage_13_out_25;
    assign stage_14_out_0 = stage_13_out_0;
    assign stage_14_out_1 = stage_13_out_1;
    assign stage_14_out_2 = stage_13_out_2;
    assign stage_14_out_3 = stage_13_out_3;
    assign stage_14_out_4 = stage_13_out_4;
    assign stage_14_out_5 = stage_13_out_5;
    assign stage_14_out_6 = stage_13_out_6;
    assign stage_14_out_7 = stage_13_out_7;
    assign stage_14_out_8 = stage_13_out_8;
    assign stage_14_out_9 = stage_13_out_9;
    assign stage_14_out_10 = stage_13_out_10;
    assign stage_14_out_12 = stage_13_out_12;
    assign stage_14_out_13 = stage_13_out_13;
    assign stage_14_out_14 = stage_13_out_14;
    assign stage_14_out_15 = stage_13_out_15;
    assign stage_14_out_16 = stage_13_out_16;
    assign stage_14_out_17 = stage_13_out_17;
    assign stage_14_out_18 = stage_13_out_18;
    assign stage_14_out_20 = stage_13_out_20;
    assign stage_14_out_22 = stage_13_out_22;
    assign stage_14_out_23 = stage_13_out_23;
    assign stage_14_out_27 = stage_13_out_27;
    assign stage_14_out_28 = stage_13_out_28;
    assign stage_14_out_32 = stage_13_out_32;
    assign stage_14_out_33 = stage_13_out_33;
    assign stage_14_out_35 = stage_13_out_35;
    assign stage_14_out_37 = stage_13_out_37;
    assign stage_14_out_38 = stage_13_out_38;
    assign stage_14_out_39 = stage_13_out_39;
    assign stage_14_out_40 = stage_13_out_40;
    assign stage_14_out_41 = stage_13_out_41;
    assign stage_14_out_42 = stage_13_out_42;
    assign stage_14_out_43 = stage_13_out_43;
    assign stage_14_out_45 = stage_13_out_45;
    assign stage_14_out_46 = stage_13_out_46;
    assign stage_14_out_47 = stage_13_out_47;
    assign stage_14_out_48 = stage_13_out_48;
    assign stage_14_out_49 = stage_13_out_49;
    assign stage_14_out_50 = stage_13_out_50;
    assign stage_14_out_51 = stage_13_out_51;
    assign stage_14_out_52 = stage_13_out_52;
    assign stage_14_out_53 = stage_13_out_53;
    assign stage_14_out_54 = stage_13_out_54;
    assign stage_14_out_55 = stage_13_out_55;
    assign stage_14_out_56 = stage_13_out_56;
    assign stage_15_out_0 = stage_14_out_0;
    assign stage_15_out_1 = stage_14_out_1;
    assign stage_15_out_2 = stage_14_out_2;
    assign stage_15_out_3 = stage_14_out_3;
    assign stage_15_out_4 = stage_14_out_4;
    assign stage_15_out_5 = stage_14_out_5;
    assign stage_15_out_6 = stage_14_out_6;
    assign stage_15_out_7 = stage_14_out_7;
    assign stage_15_out_8 = stage_14_out_8;
    assign stage_15_out_9 = stage_14_out_9;
    assign stage_15_out_10 = stage_14_out_10;
    assign stage_15_out_11 = stage_14_out_11;
    assign stage_15_out_12 = stage_14_out_12;
    assign stage_15_out_13 = stage_14_out_13;
    assign stage_15_out_14 = stage_14_out_14;
    assign stage_15_out_15 = stage_14_out_15;
    assign stage_15_out_16 = stage_14_out_16;
    assign stage_15_out_17 = stage_14_out_17;
    assign stage_15_out_18 = stage_14_out_18;
    assign stage_15_out_19 = stage_14_out_19;
    assign stage_15_out_20 = stage_14_out_20;
    assign stage_15_out_21 = stage_14_out_21;
    assign stage_15_out_22 = stage_14_out_22;
    assign stage_15_out_23 = stage_14_out_23;
    assign stage_15_out_24 = stage_14_out_24;
    assign stage_15_out_25 = stage_14_out_25;
    assign stage_15_out_26 = stage_14_out_26;
    assign stage_15_out_27 = stage_14_out_27;
    assign stage_15_out_28 = stage_14_out_28;
    assign stage_15_out_29 = stage_14_out_29;
    assign stage_15_out_30 = stage_14_out_30;
    assign stage_15_out_31 = stage_14_out_31;
    assign stage_15_out_32 = stage_14_out_32;
    assign stage_15_out_33 = stage_14_out_33;
    assign stage_15_out_34 = stage_14_out_34;
    assign stage_15_out_35 = stage_14_out_35;
    assign stage_15_out_36 = stage_14_out_36;
    assign stage_15_out_37 = stage_14_out_37;
    assign stage_15_out_38 = stage_14_out_38;
    assign stage_15_out_39 = stage_14_out_39;
    assign stage_15_out_40 = stage_14_out_40;
    assign stage_15_out_41 = stage_14_out_41;
    assign stage_15_out_42 = stage_14_out_42;
    assign stage_15_out_43 = stage_14_out_43;
    assign stage_15_out_44 = stage_14_out_44;
    assign stage_15_out_45 = stage_14_out_45;
    assign stage_15_out_46 = stage_14_out_46;
    assign stage_15_out_47 = stage_14_out_47;
    assign stage_15_out_48 = stage_14_out_48;
    assign stage_15_out_49 = stage_14_out_49;
    assign stage_15_out_50 = stage_14_out_50;
    assign stage_15_out_51 = stage_14_out_51;
    assign stage_15_out_52 = stage_14_out_52;
    assign stage_15_out_53 = stage_14_out_53;
    assign stage_15_out_54 = stage_14_out_54;
    assign stage_15_out_55 = stage_14_out_55;
    assign stage_15_out_56 = stage_14_out_56;
    assign stage_16_out_0 = stage_15_out_0;
    assign stage_16_out_1 = stage_15_out_1;
    assign stage_16_out_2 = stage_15_out_2;
    assign stage_16_out_3 = stage_15_out_3;
    assign stage_16_out_4 = stage_15_out_4;
    assign stage_16_out_5 = stage_15_out_5;
    assign stage_16_out_6 = stage_15_out_6;
    assign stage_16_out_7 = stage_15_out_7;
    assign stage_16_out_8 = stage_15_out_8;
    assign stage_16_out_9 = stage_15_out_9;
    assign stage_16_out_10 = stage_15_out_10;
    assign stage_16_out_11 = stage_15_out_11;
    assign stage_16_out_12 = stage_15_out_12;
    assign stage_16_out_13 = stage_15_out_13;
    assign stage_16_out_14 = stage_15_out_14;
    assign stage_16_out_15 = stage_15_out_15;
    assign stage_16_out_16 = stage_15_out_16;
    assign stage_16_out_17 = stage_15_out_17;
    assign stage_16_out_18 = stage_15_out_18;
    assign stage_16_out_19 = stage_15_out_19;
    assign stage_16_out_20 = stage_15_out_20;
    assign stage_16_out_21 = stage_15_out_21;
    assign stage_16_out_22 = stage_15_out_22;
    assign stage_16_out_23 = stage_15_out_23;
    assign stage_16_out_24 = stage_15_out_24;
    assign stage_16_out_25 = stage_15_out_25;
    assign stage_16_out_26 = stage_15_out_26;
    assign stage_16_out_27 = stage_15_out_27;
    assign stage_16_out_28 = stage_15_out_28;
    assign stage_16_out_29 = stage_15_out_29;
    assign stage_16_out_30 = stage_15_out_30;
    assign stage_16_out_31 = stage_15_out_31;
    assign stage_16_out_32 = stage_15_out_32;
    assign stage_16_out_33 = stage_15_out_33;
    assign stage_16_out_34 = stage_15_out_34;
    assign stage_16_out_35 = stage_15_out_35;
    assign stage_16_out_36 = stage_15_out_36;
    assign stage_16_out_37 = stage_15_out_37;
    assign stage_16_out_38 = stage_15_out_38;
    assign stage_16_out_39 = stage_15_out_39;
    assign stage_16_out_40 = stage_15_out_40;
    assign stage_16_out_41 = stage_15_out_41;
    assign stage_16_out_42 = stage_15_out_42;
    assign stage_16_out_43 = stage_15_out_43;
    assign stage_16_out_44 = stage_15_out_44;
    assign stage_16_out_45 = stage_15_out_45;
    assign stage_16_out_46 = stage_15_out_46;
    assign stage_16_out_47 = stage_15_out_47;
    assign stage_16_out_48 = stage_15_out_48;
    assign stage_16_out_49 = stage_15_out_49;
    assign stage_16_out_50 = stage_15_out_50;
    assign stage_16_out_51 = stage_15_out_51;
    assign stage_16_out_52 = stage_15_out_52;
    assign stage_16_out_53 = stage_15_out_53;
    assign stage_16_out_54 = stage_15_out_54;
    assign stage_16_out_55 = stage_15_out_55;
    assign stage_16_out_56 = stage_15_out_56;
    assign stage_17_out_0 = stage_16_out_0;
    assign stage_17_out_1 = stage_16_out_1;
    assign stage_17_out_2 = stage_16_out_2;
    assign stage_17_out_3 = stage_16_out_3;
    assign stage_17_out_4 = stage_16_out_4;
    assign stage_17_out_5 = stage_16_out_5;
    assign stage_17_out_6 = stage_16_out_6;
    assign stage_17_out_7 = stage_16_out_7;
    assign stage_17_out_8 = stage_16_out_8;
    assign stage_17_out_9 = stage_16_out_9;
    assign stage_17_out_10 = stage_16_out_10;
    assign stage_17_out_11 = stage_16_out_11;
    assign stage_17_out_12 = stage_16_out_12;
    assign stage_17_out_13 = stage_16_out_13;
    assign stage_17_out_14 = stage_16_out_14;
    assign stage_17_out_15 = stage_16_out_15;
    assign stage_17_out_16 = stage_16_out_16;
    assign stage_17_out_17 = stage_16_out_17;
    assign stage_17_out_18 = stage_16_out_18;
    assign stage_17_out_19 = stage_16_out_19;
    assign stage_17_out_20 = stage_16_out_20;
    assign stage_17_out_21 = stage_16_out_21;
    assign stage_17_out_22 = stage_16_out_22;
    assign stage_17_out_23 = stage_16_out_23;
    assign stage_17_out_24 = stage_16_out_24;
    assign stage_17_out_25 = stage_16_out_25;
    assign stage_17_out_26 = stage_16_out_26;
    assign stage_17_out_27 = stage_16_out_27;
    assign stage_17_out_28 = stage_16_out_28;
    assign stage_17_out_29 = stage_16_out_29;
    assign stage_17_out_30 = stage_16_out_30;
    assign stage_17_out_31 = stage_16_out_31;
    assign stage_17_out_32 = stage_16_out_32;
    assign stage_17_out_33 = stage_16_out_33;
    assign stage_17_out_34 = stage_16_out_34;
    assign stage_17_out_35 = stage_16_out_35;
    assign stage_17_out_36 = stage_16_out_36;
    assign stage_17_out_37 = stage_16_out_37;
    assign stage_17_out_38 = stage_16_out_38;
    assign stage_17_out_39 = stage_16_out_39;
    assign stage_17_out_40 = stage_16_out_40;
    assign stage_17_out_41 = stage_16_out_41;
    assign stage_17_out_42 = stage_16_out_42;
    assign stage_17_out_43 = stage_16_out_43;
    assign stage_17_out_44 = stage_16_out_44;
    assign stage_17_out_45 = stage_16_out_45;
    assign stage_17_out_46 = stage_16_out_46;
    assign stage_17_out_47 = stage_16_out_47;
    assign stage_17_out_48 = stage_16_out_48;
    assign stage_17_out_49 = stage_16_out_49;
    assign stage_17_out_50 = stage_16_out_50;
    assign stage_17_out_51 = stage_16_out_51;
    assign stage_17_out_52 = stage_16_out_52;
    assign stage_17_out_53 = stage_16_out_53;
    assign stage_17_out_54 = stage_16_out_54;
    assign stage_17_out_55 = stage_16_out_55;
    assign stage_17_out_56 = stage_16_out_56;
    assign stage_18_out_0 = stage_17_out_0;
    assign stage_18_out_1 = stage_17_out_1;
    assign stage_18_out_2 = stage_17_out_2;
    assign stage_18_out_3 = stage_17_out_3;
    assign stage_18_out_4 = stage_17_out_4;
    assign stage_18_out_5 = stage_17_out_5;
    assign stage_18_out_6 = stage_17_out_6;
    assign stage_18_out_7 = stage_17_out_7;
    assign stage_18_out_8 = stage_17_out_8;
    assign stage_18_out_9 = stage_17_out_9;
    assign stage_18_out_10 = stage_17_out_10;
    assign stage_18_out_11 = stage_17_out_11;
    assign stage_18_out_12 = stage_17_out_12;
    assign stage_18_out_13 = stage_17_out_13;
    assign stage_18_out_14 = stage_17_out_14;
    assign stage_18_out_15 = stage_17_out_15;
    assign stage_18_out_16 = stage_17_out_16;
    assign stage_18_out_17 = stage_17_out_17;
    assign stage_18_out_18 = stage_17_out_18;
    assign stage_18_out_19 = stage_17_out_19;
    assign stage_18_out_20 = stage_17_out_20;
    assign stage_18_out_21 = stage_17_out_21;
    assign stage_18_out_22 = stage_17_out_22;
    assign stage_18_out_23 = stage_17_out_23;
    assign stage_18_out_24 = stage_17_out_24;
    assign stage_18_out_25 = stage_17_out_25;
    assign stage_18_out_26 = stage_17_out_26;
    assign stage_18_out_27 = stage_17_out_27;
    assign stage_18_out_28 = stage_17_out_28;
    assign stage_18_out_29 = stage_17_out_29;
    assign stage_18_out_30 = stage_17_out_30;
    assign stage_18_out_31 = stage_17_out_31;
    assign stage_18_out_32 = stage_17_out_32;
    assign stage_18_out_33 = stage_17_out_33;
    assign stage_18_out_34 = stage_17_out_34;
    assign stage_18_out_35 = stage_17_out_35;
    assign stage_18_out_36 = stage_17_out_36;
    assign stage_18_out_37 = stage_17_out_37;
    assign stage_18_out_38 = stage_17_out_38;
    assign stage_18_out_39 = stage_17_out_39;
    assign stage_18_out_40 = stage_17_out_40;
    assign stage_18_out_41 = stage_17_out_41;
    assign stage_18_out_42 = stage_17_out_42;
    assign stage_18_out_43 = stage_17_out_43;
    assign stage_18_out_44 = stage_17_out_44;
    assign stage_18_out_45 = stage_17_out_45;
    assign stage_18_out_46 = stage_17_out_46;
    assign stage_18_out_47 = stage_17_out_47;
    assign stage_18_out_48 = stage_17_out_48;
    assign stage_18_out_49 = stage_17_out_49;
    assign stage_18_out_50 = stage_17_out_50;
    assign stage_18_out_51 = stage_17_out_51;
    assign stage_18_out_52 = stage_17_out_52;
    assign stage_18_out_53 = stage_17_out_53;
    assign stage_18_out_54 = stage_17_out_54;
    assign stage_18_out_55 = stage_17_out_55;
    assign stage_18_out_56 = stage_17_out_56;
    assign stage_19_out_0 = stage_18_out_0;
    assign stage_19_out_1 = stage_18_out_1;
    assign stage_19_out_2 = stage_18_out_2;
    assign stage_19_out_3 = stage_18_out_3;
    assign stage_19_out_4 = stage_18_out_4;
    assign stage_19_out_5 = stage_18_out_5;
    assign stage_19_out_6 = stage_18_out_6;
    assign stage_19_out_7 = stage_18_out_7;
    assign stage_19_out_8 = stage_18_out_8;
    assign stage_19_out_9 = stage_18_out_9;
    assign stage_19_out_10 = stage_18_out_10;
    assign stage_19_out_11 = stage_18_out_11;
    assign stage_19_out_12 = stage_18_out_12;
    assign stage_19_out_13 = stage_18_out_13;
    assign stage_19_out_14 = stage_18_out_14;
    assign stage_19_out_15 = stage_18_out_15;
    assign stage_19_out_16 = stage_18_out_16;
    assign stage_19_out_17 = stage_18_out_17;
    assign stage_19_out_18 = stage_18_out_18;
    assign stage_19_out_19 = stage_18_out_19;
    assign stage_19_out_20 = stage_18_out_20;
    assign stage_19_out_21 = stage_18_out_21;
    assign stage_19_out_22 = stage_18_out_22;
    assign stage_19_out_23 = stage_18_out_23;
    assign stage_19_out_24 = stage_18_out_24;
    assign stage_19_out_25 = stage_18_out_25;
    assign stage_19_out_26 = stage_18_out_26;
    assign stage_19_out_27 = stage_18_out_27;
    assign stage_19_out_28 = stage_18_out_28;
    assign stage_19_out_29 = stage_18_out_29;
    assign stage_19_out_30 = stage_18_out_30;
    assign stage_19_out_31 = stage_18_out_31;
    assign stage_19_out_32 = stage_18_out_32;
    assign stage_19_out_33 = stage_18_out_33;
    assign stage_19_out_34 = stage_18_out_34;
    assign stage_19_out_35 = stage_18_out_35;
    assign stage_19_out_36 = stage_18_out_36;
    assign stage_19_out_37 = stage_18_out_37;
    assign stage_19_out_38 = stage_18_out_38;
    assign stage_19_out_39 = stage_18_out_39;
    assign stage_19_out_40 = stage_18_out_40;
    assign stage_19_out_41 = stage_18_out_41;
    assign stage_19_out_42 = stage_18_out_42;
    assign stage_19_out_43 = stage_18_out_43;
    assign stage_19_out_44 = stage_18_out_44;
    assign stage_19_out_45 = stage_18_out_45;
    assign stage_19_out_46 = stage_18_out_46;
    assign stage_19_out_47 = stage_18_out_47;
    assign stage_19_out_48 = stage_18_out_48;
    assign stage_19_out_49 = stage_18_out_49;
    assign stage_19_out_50 = stage_18_out_50;
    assign stage_19_out_51 = stage_18_out_51;
    assign stage_19_out_52 = stage_18_out_52;
    assign stage_19_out_53 = stage_18_out_53;
    assign stage_19_out_54 = stage_18_out_54;
    assign stage_19_out_55 = stage_18_out_55;
    assign stage_19_out_56 = stage_18_out_56;
    assign stage_20_out_0 = stage_19_out_0;
    assign stage_20_out_1 = stage_19_out_1;
    assign stage_20_out_2 = stage_19_out_2;
    assign stage_20_out_3 = stage_19_out_3;
    assign stage_20_out_4 = stage_19_out_4;
    assign stage_20_out_5 = stage_19_out_5;
    assign stage_20_out_6 = stage_19_out_6;
    assign stage_20_out_7 = stage_19_out_7;
    assign stage_20_out_8 = stage_19_out_8;
    assign stage_20_out_9 = stage_19_out_9;
    assign stage_20_out_10 = stage_19_out_10;
    assign stage_20_out_11 = stage_19_out_11;
    assign stage_20_out_12 = stage_19_out_12;
    assign stage_20_out_13 = stage_19_out_13;
    assign stage_20_out_14 = stage_19_out_14;
    assign stage_20_out_15 = stage_19_out_15;
    assign stage_20_out_16 = stage_19_out_16;
    assign stage_20_out_17 = stage_19_out_17;
    assign stage_20_out_18 = stage_19_out_18;
    assign stage_20_out_19 = stage_19_out_19;
    assign stage_20_out_20 = stage_19_out_20;
    assign stage_20_out_21 = stage_19_out_21;
    assign stage_20_out_22 = stage_19_out_22;
    assign stage_20_out_23 = stage_19_out_23;
    assign stage_20_out_24 = stage_19_out_24;
    assign stage_20_out_25 = stage_19_out_25;
    assign stage_20_out_26 = stage_19_out_26;
    assign stage_20_out_27 = stage_19_out_27;
    assign stage_20_out_28 = stage_19_out_28;
    assign stage_20_out_29 = stage_19_out_29;
    assign stage_20_out_30 = stage_19_out_30;
    assign stage_20_out_31 = stage_19_out_31;
    assign stage_20_out_32 = stage_19_out_32;
    assign stage_20_out_33 = stage_19_out_33;
    assign stage_20_out_34 = stage_19_out_34;
    assign stage_20_out_35 = stage_19_out_35;
    assign stage_20_out_36 = stage_19_out_36;
    assign stage_20_out_37 = stage_19_out_37;
    assign stage_20_out_38 = stage_19_out_38;
    assign stage_20_out_39 = stage_19_out_39;
    assign stage_20_out_40 = stage_19_out_40;
    assign stage_20_out_41 = stage_19_out_41;
    assign stage_20_out_42 = stage_19_out_42;
    assign stage_20_out_43 = stage_19_out_43;
    assign stage_20_out_44 = stage_19_out_44;
    assign stage_20_out_45 = stage_19_out_45;
    assign stage_20_out_46 = stage_19_out_46;
    assign stage_20_out_47 = stage_19_out_47;
    assign stage_20_out_48 = stage_19_out_48;
    assign stage_20_out_49 = stage_19_out_49;
    assign stage_20_out_50 = stage_19_out_50;
    assign stage_20_out_51 = stage_19_out_51;
    assign stage_20_out_52 = stage_19_out_52;
    assign stage_20_out_53 = stage_19_out_53;
    assign stage_20_out_54 = stage_19_out_54;
    assign stage_20_out_55 = stage_19_out_55;
    assign stage_20_out_56 = stage_19_out_56;
    assign stage_21_out_0 = stage_20_out_0;
    assign stage_21_out_1 = stage_20_out_1;
    assign stage_21_out_2 = stage_20_out_2;
    assign stage_21_out_3 = stage_20_out_3;
    assign stage_21_out_4 = stage_20_out_4;
    assign stage_21_out_5 = stage_20_out_5;
    assign stage_21_out_6 = stage_20_out_6;
    assign stage_21_out_7 = stage_20_out_7;
    assign stage_21_out_8 = stage_20_out_8;
    assign stage_21_out_9 = stage_20_out_9;
    assign stage_21_out_10 = stage_20_out_10;
    assign stage_21_out_11 = stage_20_out_11;
    assign stage_21_out_12 = stage_20_out_12;
    assign stage_21_out_13 = stage_20_out_13;
    assign stage_21_out_14 = stage_20_out_14;
    assign stage_21_out_15 = stage_20_out_15;
    assign stage_21_out_16 = stage_20_out_16;
    assign stage_21_out_17 = stage_20_out_17;
    assign stage_21_out_18 = stage_20_out_18;
    assign stage_21_out_19 = stage_20_out_19;
    assign stage_21_out_20 = stage_20_out_20;
    assign stage_21_out_21 = stage_20_out_21;
    assign stage_21_out_22 = stage_20_out_22;
    assign stage_21_out_23 = stage_20_out_23;
    assign stage_21_out_24 = stage_20_out_24;
    assign stage_21_out_25 = stage_20_out_25;
    assign stage_21_out_26 = stage_20_out_26;
    assign stage_21_out_27 = stage_20_out_27;
    assign stage_21_out_28 = stage_20_out_28;
    assign stage_21_out_29 = stage_20_out_29;
    assign stage_21_out_30 = stage_20_out_30;
    assign stage_21_out_31 = stage_20_out_31;
    assign stage_21_out_32 = stage_20_out_32;
    assign stage_21_out_33 = stage_20_out_33;
    assign stage_21_out_34 = stage_20_out_34;
    assign stage_21_out_35 = stage_20_out_35;
    assign stage_21_out_36 = stage_20_out_36;
    assign stage_21_out_37 = stage_20_out_37;
    assign stage_21_out_38 = stage_20_out_38;
    assign stage_21_out_39 = stage_20_out_39;
    assign stage_21_out_40 = stage_20_out_40;
    assign stage_21_out_41 = stage_20_out_41;
    assign stage_21_out_42 = stage_20_out_42;
    assign stage_21_out_43 = stage_20_out_43;
    assign stage_21_out_44 = stage_20_out_44;
    assign stage_21_out_45 = stage_20_out_45;
    assign stage_21_out_46 = stage_20_out_46;
    assign stage_21_out_47 = stage_20_out_47;
    assign stage_21_out_48 = stage_20_out_48;
    assign stage_21_out_49 = stage_20_out_49;
    assign stage_21_out_50 = stage_20_out_50;
    assign stage_21_out_51 = stage_20_out_51;
    assign stage_21_out_52 = stage_20_out_52;
    assign stage_21_out_53 = stage_20_out_53;
    assign stage_21_out_54 = stage_20_out_54;
    assign stage_21_out_55 = stage_20_out_55;
    assign stage_21_out_56 = stage_20_out_56;
    assign stage_22_out_0 = stage_21_out_0;
    assign stage_22_out_1 = stage_21_out_1;
    assign stage_22_out_2 = stage_21_out_2;
    assign stage_22_out_3 = stage_21_out_3;
    assign stage_22_out_4 = stage_21_out_4;
    assign stage_22_out_5 = stage_21_out_5;
    assign stage_22_out_6 = stage_21_out_6;
    assign stage_22_out_7 = stage_21_out_7;
    assign stage_22_out_8 = stage_21_out_8;
    assign stage_22_out_9 = stage_21_out_9;
    assign stage_22_out_10 = stage_21_out_10;
    assign stage_22_out_11 = stage_21_out_11;
    assign stage_22_out_12 = stage_21_out_12;
    assign stage_22_out_13 = stage_21_out_13;
    assign stage_22_out_14 = stage_21_out_14;
    assign stage_22_out_15 = stage_21_out_15;
    assign stage_22_out_16 = stage_21_out_16;
    assign stage_22_out_17 = stage_21_out_17;
    assign stage_22_out_18 = stage_21_out_18;
    assign stage_22_out_19 = stage_21_out_19;
    assign stage_22_out_20 = stage_21_out_20;
    assign stage_22_out_21 = stage_21_out_21;
    assign stage_22_out_22 = stage_21_out_22;
    assign stage_22_out_23 = stage_21_out_23;
    assign stage_22_out_24 = stage_21_out_24;
    assign stage_22_out_25 = stage_21_out_25;
    assign stage_22_out_26 = stage_21_out_26;
    assign stage_22_out_27 = stage_21_out_27;
    assign stage_22_out_28 = stage_21_out_28;
    assign stage_22_out_29 = stage_21_out_29;
    assign stage_22_out_30 = stage_21_out_30;
    assign stage_22_out_31 = stage_21_out_31;
    assign stage_22_out_32 = stage_21_out_32;
    assign stage_22_out_33 = stage_21_out_33;
    assign stage_22_out_34 = stage_21_out_34;
    assign stage_22_out_35 = stage_21_out_35;
    assign stage_22_out_36 = stage_21_out_36;
    assign stage_22_out_37 = stage_21_out_37;
    assign stage_22_out_38 = stage_21_out_38;
    assign stage_22_out_39 = stage_21_out_39;
    assign stage_22_out_40 = stage_21_out_40;
    assign stage_22_out_41 = stage_21_out_41;
    assign stage_22_out_42 = stage_21_out_42;
    assign stage_22_out_43 = stage_21_out_43;
    assign stage_22_out_44 = stage_21_out_44;
    assign stage_22_out_45 = stage_21_out_45;
    assign stage_22_out_46 = stage_21_out_46;
    assign stage_22_out_47 = stage_21_out_47;
    assign stage_22_out_48 = stage_21_out_48;
    assign stage_22_out_49 = stage_21_out_49;
    assign stage_22_out_50 = stage_21_out_50;
    assign stage_22_out_51 = stage_21_out_51;
    assign stage_22_out_52 = stage_21_out_52;
    assign stage_22_out_53 = stage_21_out_53;
    assign stage_22_out_54 = stage_21_out_54;
    assign stage_22_out_55 = stage_21_out_55;
    assign stage_22_out_56 = stage_21_out_56;
    assign stage_23_out_0 = stage_22_out_0;
    assign stage_23_out_1 = stage_22_out_1;
    assign stage_23_out_2 = stage_22_out_2;
    assign stage_23_out_3 = stage_22_out_3;
    assign stage_23_out_4 = stage_22_out_4;
    assign stage_23_out_5 = stage_22_out_5;
    assign stage_23_out_6 = stage_22_out_6;
    assign stage_23_out_7 = stage_22_out_7;
    assign stage_23_out_8 = stage_22_out_8;
    assign stage_23_out_9 = stage_22_out_9;
    assign stage_23_out_10 = stage_22_out_10;
    assign stage_23_out_11 = stage_22_out_11;
    assign stage_23_out_12 = stage_22_out_12;
    assign stage_23_out_13 = stage_22_out_13;
    assign stage_23_out_14 = stage_22_out_14;
    assign stage_23_out_15 = stage_22_out_15;
    assign stage_23_out_16 = stage_22_out_16;
    assign stage_23_out_17 = stage_22_out_17;
    assign stage_23_out_18 = stage_22_out_18;
    assign stage_23_out_19 = stage_22_out_19;
    assign stage_23_out_20 = stage_22_out_20;
    assign stage_23_out_21 = stage_22_out_21;
    assign stage_23_out_22 = stage_22_out_22;
    assign stage_23_out_23 = stage_22_out_23;
    assign stage_23_out_24 = stage_22_out_24;
    assign stage_23_out_25 = stage_22_out_25;
    assign stage_23_out_26 = stage_22_out_26;
    assign stage_23_out_27 = stage_22_out_27;
    assign stage_23_out_28 = stage_22_out_28;
    assign stage_23_out_29 = stage_22_out_29;
    assign stage_23_out_30 = stage_22_out_30;
    assign stage_23_out_31 = stage_22_out_31;
    assign stage_23_out_32 = stage_22_out_32;
    assign stage_23_out_33 = stage_22_out_33;
    assign stage_23_out_34 = stage_22_out_34;
    assign stage_23_out_35 = stage_22_out_35;
    assign stage_23_out_36 = stage_22_out_36;
    assign stage_23_out_37 = stage_22_out_37;
    assign stage_23_out_38 = stage_22_out_38;
    assign stage_23_out_39 = stage_22_out_39;
    assign stage_23_out_40 = stage_22_out_40;
    assign stage_23_out_41 = stage_22_out_41;
    assign stage_23_out_42 = stage_22_out_42;
    assign stage_23_out_43 = stage_22_out_43;
    assign stage_23_out_44 = stage_22_out_44;
    assign stage_23_out_45 = stage_22_out_45;
    assign stage_23_out_46 = stage_22_out_46;
    assign stage_23_out_47 = stage_22_out_47;
    assign stage_23_out_48 = stage_22_out_48;
    assign stage_23_out_49 = stage_22_out_49;
    assign stage_23_out_50 = stage_22_out_50;
    assign stage_23_out_51 = stage_22_out_51;
    assign stage_23_out_52 = stage_22_out_52;
    assign stage_23_out_53 = stage_22_out_53;
    assign stage_23_out_54 = stage_22_out_54;
    assign stage_23_out_55 = stage_22_out_55;
    assign stage_23_out_56 = stage_22_out_56;
    assign stage_24_out_0 = stage_23_out_0;
    assign stage_24_out_1 = stage_23_out_1;
    assign stage_24_out_2 = stage_23_out_2;
    assign stage_24_out_3 = stage_23_out_3;
    assign stage_24_out_4 = stage_23_out_4;
    assign stage_24_out_5 = stage_23_out_5;
    assign stage_24_out_6 = stage_23_out_6;
    assign stage_24_out_7 = stage_23_out_7;
    assign stage_24_out_8 = stage_23_out_8;
    assign stage_24_out_9 = stage_23_out_9;
    assign stage_24_out_10 = stage_23_out_10;
    assign stage_24_out_11 = stage_23_out_11;
    assign stage_24_out_12 = stage_23_out_12;
    assign stage_24_out_13 = stage_23_out_13;
    assign stage_24_out_14 = stage_23_out_14;
    assign stage_24_out_15 = stage_23_out_15;
    assign stage_24_out_16 = stage_23_out_16;
    assign stage_24_out_17 = stage_23_out_17;
    assign stage_24_out_18 = stage_23_out_18;
    assign stage_24_out_19 = stage_23_out_19;
    assign stage_24_out_20 = stage_23_out_20;
    assign stage_24_out_21 = stage_23_out_21;
    assign stage_24_out_22 = stage_23_out_22;
    assign stage_24_out_23 = stage_23_out_23;
    assign stage_24_out_24 = stage_23_out_24;
    assign stage_24_out_25 = stage_23_out_25;
    assign stage_24_out_26 = stage_23_out_26;
    assign stage_24_out_27 = stage_23_out_27;
    assign stage_24_out_28 = stage_23_out_28;
    assign stage_24_out_29 = stage_23_out_29;
    assign stage_24_out_30 = stage_23_out_30;
    assign stage_24_out_31 = stage_23_out_31;
    assign stage_24_out_32 = stage_23_out_32;
    assign stage_24_out_33 = stage_23_out_33;
    assign stage_24_out_34 = stage_23_out_34;
    assign stage_24_out_35 = stage_23_out_35;
    assign stage_24_out_36 = stage_23_out_36;
    assign stage_24_out_37 = stage_23_out_37;
    assign stage_24_out_38 = stage_23_out_38;
    assign stage_24_out_39 = stage_23_out_39;
    assign stage_24_out_40 = stage_23_out_40;
    assign stage_24_out_41 = stage_23_out_41;
    assign stage_24_out_42 = stage_23_out_42;
    assign stage_24_out_43 = stage_23_out_43;
    assign stage_24_out_44 = stage_23_out_44;
    assign stage_24_out_45 = stage_23_out_45;
    assign stage_24_out_46 = stage_23_out_46;
    assign stage_24_out_47 = stage_23_out_47;
    assign stage_24_out_48 = stage_23_out_48;
    assign stage_24_out_49 = stage_23_out_49;
    assign stage_24_out_50 = stage_23_out_50;
    assign stage_24_out_51 = stage_23_out_51;
    assign stage_24_out_52 = stage_23_out_52;
    assign stage_24_out_53 = stage_23_out_53;
    assign stage_24_out_54 = stage_23_out_54;
    assign stage_24_out_55 = stage_23_out_55;
    assign stage_24_out_56 = stage_23_out_56;
    assign stage_25_out_0 = stage_24_out_0;
    assign stage_25_out_1 = stage_24_out_1;
    assign stage_25_out_2 = stage_24_out_2;
    assign stage_25_out_3 = stage_24_out_3;
    assign stage_25_out_4 = stage_24_out_4;
    assign stage_25_out_5 = stage_24_out_5;
    assign stage_25_out_6 = stage_24_out_6;
    assign stage_25_out_7 = stage_24_out_7;
    assign stage_25_out_8 = stage_24_out_8;
    assign stage_25_out_9 = stage_24_out_9;
    assign stage_25_out_10 = stage_24_out_10;
    assign stage_25_out_11 = stage_24_out_11;
    assign stage_25_out_12 = stage_24_out_12;
    assign stage_25_out_13 = stage_24_out_13;
    assign stage_25_out_14 = stage_24_out_14;
    assign stage_25_out_15 = stage_24_out_15;
    assign stage_25_out_16 = stage_24_out_16;
    assign stage_25_out_17 = stage_24_out_17;
    assign stage_25_out_18 = stage_24_out_18;
    assign stage_25_out_19 = stage_24_out_19;
    assign stage_25_out_20 = stage_24_out_20;
    assign stage_25_out_21 = stage_24_out_21;
    assign stage_25_out_22 = stage_24_out_22;
    assign stage_25_out_23 = stage_24_out_23;
    assign stage_25_out_24 = stage_24_out_24;
    assign stage_25_out_25 = stage_24_out_25;
    assign stage_25_out_26 = stage_24_out_26;
    assign stage_25_out_27 = stage_24_out_27;
    assign stage_25_out_28 = stage_24_out_28;
    assign stage_25_out_29 = stage_24_out_29;
    assign stage_25_out_30 = stage_24_out_30;
    assign stage_25_out_31 = stage_24_out_31;
    assign stage_25_out_32 = stage_24_out_32;
    assign stage_25_out_33 = stage_24_out_33;
    assign stage_25_out_34 = stage_24_out_34;
    assign stage_25_out_35 = stage_24_out_35;
    assign stage_25_out_36 = stage_24_out_36;
    assign stage_25_out_37 = stage_24_out_37;
    assign stage_25_out_38 = stage_24_out_38;
    assign stage_25_out_39 = stage_24_out_39;
    assign stage_25_out_40 = stage_24_out_40;
    assign stage_25_out_41 = stage_24_out_41;
    assign stage_25_out_42 = stage_24_out_42;
    assign stage_25_out_43 = stage_24_out_43;
    assign stage_25_out_44 = stage_24_out_44;
    assign stage_25_out_45 = stage_24_out_45;
    assign stage_25_out_46 = stage_24_out_46;
    assign stage_25_out_47 = stage_24_out_47;
    assign stage_25_out_48 = stage_24_out_48;
    assign stage_25_out_49 = stage_24_out_49;
    assign stage_25_out_50 = stage_24_out_50;
    assign stage_25_out_51 = stage_24_out_51;
    assign stage_25_out_52 = stage_24_out_52;
    assign stage_25_out_53 = stage_24_out_53;
    assign stage_25_out_54 = stage_24_out_54;
    assign stage_25_out_55 = stage_24_out_55;
    assign stage_25_out_56 = stage_24_out_56;
    assign sort_0 = stage_25_out_0;
    assign sort_1 = stage_25_out_1;
    assign sort_2 = stage_25_out_2;
    assign sort_3 = stage_25_out_3;
    assign sort_4 = stage_25_out_4;
    assign sort_5 = stage_25_out_5;
    assign sort_6 = stage_25_out_6;
    assign sort_7 = stage_25_out_7;
    assign sort_8 = stage_25_out_8;
    assign sort_9 = stage_25_out_9;
    assign sort_10 = stage_25_out_10;
    assign sort_11 = stage_25_out_11;
    assign sort_12 = stage_25_out_12;
    assign sort_13 = stage_25_out_13;
    assign sort_14 = stage_25_out_14;
    assign sort_15 = stage_25_out_15;
    assign sort_16 = stage_25_out_16;
    assign sort_17 = stage_25_out_17;
    assign sort_18 = stage_25_out_18;
    assign sort_19 = stage_25_out_19;
    assign sort_20 = stage_25_out_20;
    assign sort_21 = stage_25_out_21;
    assign sort_22 = stage_25_out_22;
    assign sort_23 = stage_25_out_23;
    assign sort_24 = stage_25_out_24;
    assign sort_25 = stage_25_out_25;
    assign sort_26 = stage_25_out_26;
    assign sort_27 = stage_25_out_27;
    assign sort_28 = stage_25_out_28;
    assign sort_29 = stage_25_out_29;
    assign sort_30 = stage_25_out_30;
    assign sort_31 = stage_25_out_31;
    assign sort_32 = stage_25_out_32;
    assign sort_33 = stage_25_out_33;
    assign sort_34 = stage_25_out_34;
    assign sort_35 = stage_25_out_35;
    assign sort_36 = stage_25_out_36;
    assign sort_37 = stage_25_out_37;
    assign sort_38 = stage_25_out_38;
    assign sort_39 = stage_25_out_39;
    assign sort_40 = stage_25_out_40;
    assign sort_41 = stage_25_out_41;
    assign sort_42 = stage_25_out_42;
    assign sort_43 = stage_25_out_43;
    assign sort_44 = stage_25_out_44;
    assign sort_45 = stage_25_out_45;
    assign sort_46 = stage_25_out_46;
    assign sort_47 = stage_25_out_47;
    assign sort_48 = stage_25_out_48;
    assign sort_49 = stage_25_out_49;
    assign sort_50 = stage_25_out_50;
    assign sort_51 = stage_25_out_51;
    assign sort_52 = stage_25_out_52;
    assign sort_53 = stage_25_out_53;
    assign sort_54 = stage_25_out_54;
    assign sort_55 = stage_25_out_55;
    assign sort_56 = stage_25_out_56;
endmodule

module median_57_292_26_tb;

    logic clk;
    data_t data_0;
    data_t data_1;
    data_t data_2;
    data_t data_3;
    data_t data_4;
    data_t data_5;
    data_t data_6;
    data_t data_7;
    data_t data_8;
    data_t data_9;
    data_t data_10;
    data_t data_11;
    data_t data_12;
    data_t data_13;
    data_t data_14;
    data_t data_15;
    data_t data_16;
    data_t data_17;
    data_t data_18;
    data_t data_19;
    data_t data_20;
    data_t data_21;
    data_t data_22;
    data_t data_23;
    data_t data_24;
    data_t data_25;
    data_t data_26;
    data_t data_27;
    data_t data_28;
    data_t data_29;
    data_t data_30;
    data_t data_31;
    data_t data_32;
    data_t data_33;
    data_t data_34;
    data_t data_35;
    data_t data_36;
    data_t data_37;
    data_t data_38;
    data_t data_39;
    data_t data_40;
    data_t data_41;
    data_t data_42;
    data_t data_43;
    data_t data_44;
    data_t data_45;
    data_t data_46;
    data_t data_47;
    data_t data_48;
    data_t data_49;
    data_t data_50;
    data_t data_51;
    data_t data_52;
    data_t data_53;
    data_t data_54;
    data_t data_55;
    data_t data_56;
    data_t sort_0;
    data_t sort_1;
    data_t sort_2;
    data_t sort_3;
    data_t sort_4;
    data_t sort_5;
    data_t sort_6;
    data_t sort_7;
    data_t sort_8;
    data_t sort_9;
    data_t sort_10;
    data_t sort_11;
    data_t sort_12;
    data_t sort_13;
    data_t sort_14;
    data_t sort_15;
    data_t sort_16;
    data_t sort_17;
    data_t sort_18;
    data_t sort_19;
    data_t sort_20;
    data_t sort_21;
    data_t sort_22;
    data_t sort_23;
    data_t sort_24;
    data_t sort_25;
    data_t sort_26;
    data_t sort_27;
    data_t sort_28;
    data_t sort_29;
    data_t sort_30;
    data_t sort_31;
    data_t sort_32;
    data_t sort_33;
    data_t sort_34;
    data_t sort_35;
    data_t sort_36;
    data_t sort_37;
    data_t sort_38;
    data_t sort_39;
    data_t sort_40;
    data_t sort_41;
    data_t sort_42;
    data_t sort_43;
    data_t sort_44;
    data_t sort_45;
    data_t sort_46;
    data_t sort_47;
    data_t sort_48;
    data_t sort_49;
    data_t sort_50;
    data_t sort_51;
    data_t sort_52;
    data_t sort_53;
    data_t sort_54;
    data_t sort_55;
    data_t sort_56;

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Instantiate DUT
    median_57_292_26 dut (
        .clk(clk),
        .data_0(data_0),
        .data_1(data_1),
        .data_2(data_2),
        .data_3(data_3),
        .data_4(data_4),
        .data_5(data_5),
        .data_6(data_6),
        .data_7(data_7),
        .data_8(data_8),
        .data_9(data_9),
        .data_10(data_10),
        .data_11(data_11),
        .data_12(data_12),
        .data_13(data_13),
        .data_14(data_14),
        .data_15(data_15),
        .data_16(data_16),
        .data_17(data_17),
        .data_18(data_18),
        .data_19(data_19),
        .data_20(data_20),
        .data_21(data_21),
        .data_22(data_22),
        .data_23(data_23),
        .data_24(data_24),
        .data_25(data_25),
        .data_26(data_26),
        .data_27(data_27),
        .data_28(data_28),
        .data_29(data_29),
        .data_30(data_30),
        .data_31(data_31),
        .data_32(data_32),
        .data_33(data_33),
        .data_34(data_34),
        .data_35(data_35),
        .data_36(data_36),
        .data_37(data_37),
        .data_38(data_38),
        .data_39(data_39),
        .data_40(data_40),
        .data_41(data_41),
        .data_42(data_42),
        .data_43(data_43),
        .data_44(data_44),
        .data_45(data_45),
        .data_46(data_46),
        .data_47(data_47),
        .data_48(data_48),
        .data_49(data_49),
        .data_50(data_50),
        .data_51(data_51),
        .data_52(data_52),
        .data_53(data_53),
        .data_54(data_54),
        .data_55(data_55),
        .data_56(data_56),
        .sort_0(sort_0),
        .sort_1(sort_1),
        .sort_2(sort_2),
        .sort_3(sort_3),
        .sort_4(sort_4),
        .sort_5(sort_5),
        .sort_6(sort_6),
        .sort_7(sort_7),
        .sort_8(sort_8),
        .sort_9(sort_9),
        .sort_10(sort_10),
        .sort_11(sort_11),
        .sort_12(sort_12),
        .sort_13(sort_13),
        .sort_14(sort_14),
        .sort_15(sort_15),
        .sort_16(sort_16),
        .sort_17(sort_17),
        .sort_18(sort_18),
        .sort_19(sort_19),
        .sort_20(sort_20),
        .sort_21(sort_21),
        .sort_22(sort_22),
        .sort_23(sort_23),
        .sort_24(sort_24),
        .sort_25(sort_25),
        .sort_26(sort_26),
        .sort_27(sort_27),
        .sort_28(sort_28),
        .sort_29(sort_29),
        .sort_30(sort_30),
        .sort_31(sort_31),
        .sort_32(sort_32),
        .sort_33(sort_33),
        .sort_34(sort_34),
        .sort_35(sort_35),
        .sort_36(sort_36),
        .sort_37(sort_37),
        .sort_38(sort_38),
        .sort_39(sort_39),
        .sort_40(sort_40),
        .sort_41(sort_41),
        .sort_42(sort_42),
        .sort_43(sort_43),
        .sort_44(sort_44),
        .sort_45(sort_45),
        .sort_46(sort_46),
        .sort_47(sort_47),
        .sort_48(sort_48),
        .sort_49(sort_49),
        .sort_50(sort_50),
        .sort_51(sort_51),
        .sort_52(sort_52),
        .sort_53(sort_53),
        .sort_54(sort_54),
        .sort_55(sort_55),
        .sort_56(sort_56)
    );

    // Apply random inputs
    initial begin
        repeat (100) begin
            @(posedge clk);
            data_0 = $urandom;
            data_1 = $urandom;
            data_2 = $urandom;
            data_3 = $urandom;
            data_4 = $urandom;
            data_5 = $urandom;
            data_6 = $urandom;
            data_7 = $urandom;
            data_8 = $urandom;
            data_9 = $urandom;
            data_10 = $urandom;
            data_11 = $urandom;
            data_12 = $urandom;
            data_13 = $urandom;
            data_14 = $urandom;
            data_15 = $urandom;
            data_16 = $urandom;
            data_17 = $urandom;
            data_18 = $urandom;
            data_19 = $urandom;
            data_20 = $urandom;
            data_21 = $urandom;
            data_22 = $urandom;
            data_23 = $urandom;
            data_24 = $urandom;
            data_25 = $urandom;
            data_26 = $urandom;
            data_27 = $urandom;
            data_28 = $urandom;
            data_29 = $urandom;
            data_30 = $urandom;
            data_31 = $urandom;
            data_32 = $urandom;
            data_33 = $urandom;
            data_34 = $urandom;
            data_35 = $urandom;
            data_36 = $urandom;
            data_37 = $urandom;
            data_38 = $urandom;
            data_39 = $urandom;
            data_40 = $urandom;
            data_41 = $urandom;
            data_42 = $urandom;
            data_43 = $urandom;
            data_44 = $urandom;
            data_45 = $urandom;
            data_46 = $urandom;
            data_47 = $urandom;
            data_48 = $urandom;
            data_49 = $urandom;
            data_50 = $urandom;
            data_51 = $urandom;
            data_52 = $urandom;
            data_53 = $urandom;
            data_54 = $urandom;
            data_55 = $urandom;
            data_56 = $urandom;
        end
        #100 $finish;
    end

    // Verification logic
    localparam int latency = 0;
    integer cycle_count = 0;
    integer success_count = 0;
    integer failure_count = 0;
    always @(posedge clk) begin
        cycle_count <= cycle_count + 1;
        if (cycle_count > latency) begin
            if (sort_0 <= sort_1 && sort_1 <= sort_2 && sort_2 <= sort_3 && sort_3 <= sort_4 && sort_4 <= sort_5 && sort_5 <= sort_6 && sort_6 <= sort_7 && sort_7 <= sort_8 && sort_8 <= sort_9 && sort_9 <= sort_10 && sort_10 <= sort_11 && sort_11 <= sort_12 && sort_12 <= sort_13 && sort_13 <= sort_14 && sort_14 <= sort_15 && sort_15 <= sort_16 && sort_16 <= sort_17 && sort_17 <= sort_18 && sort_18 <= sort_19 && sort_19 <= sort_20 && sort_20 <= sort_21 && sort_21 <= sort_22 && sort_22 <= sort_23 && sort_23 <= sort_24 && sort_24 <= sort_25 && sort_25 <= sort_26 && sort_26 <= sort_27 && sort_27 <= sort_28 && sort_28 <= sort_29 && sort_29 <= sort_30 && sort_30 <= sort_31 && sort_31 <= sort_32 && sort_32 <= sort_33 && sort_33 <= sort_34 && sort_34 <= sort_35 && sort_35 <= sort_36 && sort_36 <= sort_37 && sort_37 <= sort_38 && sort_38 <= sort_39 && sort_39 <= sort_40 && sort_40 <= sort_41 && sort_41 <= sort_42 && sort_42 <= sort_43 && sort_43 <= sort_44 && sort_44 <= sort_45 && sort_45 <= sort_46 && sort_46 <= sort_47 && sort_47 <= sort_48 && sort_48 <= sort_49 && sort_49 <= sort_50 && sort_50 <= sort_51 && sort_51 <= sort_52 && sort_52 <= sort_53 && sort_53 <= sort_54 && sort_54 <= sort_55 && sort_55 <= sort_56) begin
                success_count <= success_count + 1;
            end else begin
                failure_count <= failure_count + 1;
            end
            $display("Cycle: %0d, Success: %0d, Failure: %0d", cycle_count, success_count, failure_count);
        end
    end

endmodule