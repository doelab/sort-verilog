typedef logic [31:0] data_t;

module sort_34_209_17 (
    input logic clk,
    input data_t data_0,
    input data_t data_1,
    input data_t data_2,
    input data_t data_3,
    input data_t data_4,
    input data_t data_5,
    input data_t data_6,
    input data_t data_7,
    input data_t data_8,
    input data_t data_9,
    input data_t data_10,
    input data_t data_11,
    input data_t data_12,
    input data_t data_13,
    input data_t data_14,
    input data_t data_15,
    input data_t data_16,
    input data_t data_17,
    input data_t data_18,
    input data_t data_19,
    input data_t data_20,
    input data_t data_21,
    input data_t data_22,
    input data_t data_23,
    input data_t data_24,
    input data_t data_25,
    input data_t data_26,
    input data_t data_27,
    input data_t data_28,
    input data_t data_29,
    input data_t data_30,
    input data_t data_31,
    input data_t data_32,
    input data_t data_33,
    output data_t sort_0,
    output data_t sort_1,
    output data_t sort_2,
    output data_t sort_3,
    output data_t sort_4,
    output data_t sort_5,
    output data_t sort_6,
    output data_t sort_7,
    output data_t sort_8,
    output data_t sort_9,
    output data_t sort_10,
    output data_t sort_11,
    output data_t sort_12,
    output data_t sort_13,
    output data_t sort_14,
    output data_t sort_15,
    output data_t sort_16,
    output data_t sort_17,
    output data_t sort_18,
    output data_t sort_19,
    output data_t sort_20,
    output data_t sort_21,
    output data_t sort_22,
    output data_t sort_23,
    output data_t sort_24,
    output data_t sort_25,
    output data_t sort_26,
    output data_t sort_27,
    output data_t sort_28,
    output data_t sort_29,
    output data_t sort_30,
    output data_t sort_31,
    output data_t sort_32,
    output data_t sort_33
);

     logic [31:0] stage_0_out_0;
     logic [31:0] stage_0_out_1;
     logic [31:0] stage_0_out_2;
     logic [31:0] stage_0_out_3;
     logic [31:0] stage_0_out_4;
     logic [31:0] stage_0_out_5;
     logic [31:0] stage_0_out_6;
     logic [31:0] stage_0_out_7;
     logic [31:0] stage_0_out_8;
     logic [31:0] stage_0_out_9;
     logic [31:0] stage_0_out_10;
     logic [31:0] stage_0_out_11;
     logic [31:0] stage_0_out_12;
     logic [31:0] stage_0_out_13;
     logic [31:0] stage_0_out_14;
     logic [31:0] stage_0_out_15;
     logic [31:0] stage_0_out_16;
     logic [31:0] stage_0_out_17;
     logic [31:0] stage_0_out_18;
     logic [31:0] stage_0_out_19;
     logic [31:0] stage_0_out_20;
     logic [31:0] stage_0_out_21;
     logic [31:0] stage_0_out_22;
     logic [31:0] stage_0_out_23;
     logic [31:0] stage_0_out_24;
     logic [31:0] stage_0_out_25;
     logic [31:0] stage_0_out_26;
     logic [31:0] stage_0_out_27;
     logic [31:0] stage_0_out_28;
     logic [31:0] stage_0_out_29;
     logic [31:0] stage_0_out_30;
     logic [31:0] stage_0_out_31;
     logic [31:0] stage_0_out_32;
     logic [31:0] stage_0_out_33;
     logic [31:0] stage_1_out_0;
     logic [31:0] stage_1_out_1;
     logic [31:0] stage_1_out_2;
     logic [31:0] stage_1_out_3;
     logic [31:0] stage_1_out_4;
     logic [31:0] stage_1_out_5;
     logic [31:0] stage_1_out_6;
     logic [31:0] stage_1_out_7;
     logic [31:0] stage_1_out_8;
     logic [31:0] stage_1_out_9;
     logic [31:0] stage_1_out_10;
     logic [31:0] stage_1_out_11;
     logic [31:0] stage_1_out_12;
     logic [31:0] stage_1_out_13;
     logic [31:0] stage_1_out_14;
     logic [31:0] stage_1_out_15;
     logic [31:0] stage_1_out_16;
     logic [31:0] stage_1_out_17;
     logic [31:0] stage_1_out_18;
     logic [31:0] stage_1_out_19;
     logic [31:0] stage_1_out_20;
     logic [31:0] stage_1_out_21;
     logic [31:0] stage_1_out_22;
     logic [31:0] stage_1_out_23;
     logic [31:0] stage_1_out_24;
     logic [31:0] stage_1_out_25;
     logic [31:0] stage_1_out_26;
     logic [31:0] stage_1_out_27;
     logic [31:0] stage_1_out_28;
     logic [31:0] stage_1_out_29;
     logic [31:0] stage_1_out_30;
     logic [31:0] stage_1_out_31;
     logic [31:0] stage_1_out_32;
     logic [31:0] stage_1_out_33;
     logic [31:0] stage_2_out_0;
     logic [31:0] stage_2_out_1;
     logic [31:0] stage_2_out_2;
     logic [31:0] stage_2_out_3;
     logic [31:0] stage_2_out_4;
     logic [31:0] stage_2_out_5;
     logic [31:0] stage_2_out_6;
     logic [31:0] stage_2_out_7;
     logic [31:0] stage_2_out_8;
     logic [31:0] stage_2_out_9;
     logic [31:0] stage_2_out_10;
     logic [31:0] stage_2_out_11;
     logic [31:0] stage_2_out_12;
     logic [31:0] stage_2_out_13;
     logic [31:0] stage_2_out_14;
     logic [31:0] stage_2_out_15;
     logic [31:0] stage_2_out_16;
     logic [31:0] stage_2_out_17;
     logic [31:0] stage_2_out_18;
     logic [31:0] stage_2_out_19;
     logic [31:0] stage_2_out_20;
     logic [31:0] stage_2_out_21;
     logic [31:0] stage_2_out_22;
     logic [31:0] stage_2_out_23;
     logic [31:0] stage_2_out_24;
     logic [31:0] stage_2_out_25;
     logic [31:0] stage_2_out_26;
     logic [31:0] stage_2_out_27;
     logic [31:0] stage_2_out_28;
     logic [31:0] stage_2_out_29;
     logic [31:0] stage_2_out_30;
     logic [31:0] stage_2_out_31;
     logic [31:0] stage_2_out_32;
     logic [31:0] stage_2_out_33;
     logic [31:0] stage_3_out_0;
     logic [31:0] stage_3_out_1;
     logic [31:0] stage_3_out_2;
     logic [31:0] stage_3_out_3;
     logic [31:0] stage_3_out_4;
     logic [31:0] stage_3_out_5;
     logic [31:0] stage_3_out_6;
     logic [31:0] stage_3_out_7;
     logic [31:0] stage_3_out_8;
     logic [31:0] stage_3_out_9;
     logic [31:0] stage_3_out_10;
     logic [31:0] stage_3_out_11;
     logic [31:0] stage_3_out_12;
     logic [31:0] stage_3_out_13;
     logic [31:0] stage_3_out_14;
     logic [31:0] stage_3_out_15;
     logic [31:0] stage_3_out_16;
     logic [31:0] stage_3_out_17;
     logic [31:0] stage_3_out_18;
     logic [31:0] stage_3_out_19;
     logic [31:0] stage_3_out_20;
     logic [31:0] stage_3_out_21;
     logic [31:0] stage_3_out_22;
     logic [31:0] stage_3_out_23;
     logic [31:0] stage_3_out_24;
     logic [31:0] stage_3_out_25;
     logic [31:0] stage_3_out_26;
     logic [31:0] stage_3_out_27;
     logic [31:0] stage_3_out_28;
     logic [31:0] stage_3_out_29;
     logic [31:0] stage_3_out_30;
     logic [31:0] stage_3_out_31;
     logic [31:0] stage_3_out_32;
     logic [31:0] stage_3_out_33;
     logic [31:0] stage_4_out_0;
     logic [31:0] stage_4_out_1;
     logic [31:0] stage_4_out_2;
     logic [31:0] stage_4_out_3;
     logic [31:0] stage_4_out_4;
     logic [31:0] stage_4_out_5;
     logic [31:0] stage_4_out_6;
     logic [31:0] stage_4_out_7;
     logic [31:0] stage_4_out_8;
     logic [31:0] stage_4_out_9;
     logic [31:0] stage_4_out_10;
     logic [31:0] stage_4_out_11;
     logic [31:0] stage_4_out_12;
     logic [31:0] stage_4_out_13;
     logic [31:0] stage_4_out_14;
     logic [31:0] stage_4_out_15;
     logic [31:0] stage_4_out_16;
     logic [31:0] stage_4_out_17;
     logic [31:0] stage_4_out_18;
     logic [31:0] stage_4_out_19;
     logic [31:0] stage_4_out_20;
     logic [31:0] stage_4_out_21;
     logic [31:0] stage_4_out_22;
     logic [31:0] stage_4_out_23;
     logic [31:0] stage_4_out_24;
     logic [31:0] stage_4_out_25;
     logic [31:0] stage_4_out_26;
     logic [31:0] stage_4_out_27;
     logic [31:0] stage_4_out_28;
     logic [31:0] stage_4_out_29;
     logic [31:0] stage_4_out_30;
     logic [31:0] stage_4_out_31;
     logic [31:0] stage_4_out_32;
     logic [31:0] stage_4_out_33;
     logic [31:0] stage_5_out_0;
     logic [31:0] stage_5_out_1;
     logic [31:0] stage_5_out_2;
     logic [31:0] stage_5_out_3;
     logic [31:0] stage_5_out_4;
     logic [31:0] stage_5_out_5;
     logic [31:0] stage_5_out_6;
     logic [31:0] stage_5_out_7;
     logic [31:0] stage_5_out_8;
     logic [31:0] stage_5_out_9;
     logic [31:0] stage_5_out_10;
     logic [31:0] stage_5_out_11;
     logic [31:0] stage_5_out_12;
     logic [31:0] stage_5_out_13;
     logic [31:0] stage_5_out_14;
     logic [31:0] stage_5_out_15;
     logic [31:0] stage_5_out_16;
     logic [31:0] stage_5_out_17;
     logic [31:0] stage_5_out_18;
     logic [31:0] stage_5_out_19;
     logic [31:0] stage_5_out_20;
     logic [31:0] stage_5_out_21;
     logic [31:0] stage_5_out_22;
     logic [31:0] stage_5_out_23;
     logic [31:0] stage_5_out_24;
     logic [31:0] stage_5_out_25;
     logic [31:0] stage_5_out_26;
     logic [31:0] stage_5_out_27;
     logic [31:0] stage_5_out_28;
     logic [31:0] stage_5_out_29;
     logic [31:0] stage_5_out_30;
     logic [31:0] stage_5_out_31;
     logic [31:0] stage_5_out_32;
     logic [31:0] stage_5_out_33;
     logic [31:0] stage_6_out_0;
     logic [31:0] stage_6_out_1;
     logic [31:0] stage_6_out_2;
     logic [31:0] stage_6_out_3;
     logic [31:0] stage_6_out_4;
     logic [31:0] stage_6_out_5;
     logic [31:0] stage_6_out_6;
     logic [31:0] stage_6_out_7;
     logic [31:0] stage_6_out_8;
     logic [31:0] stage_6_out_9;
     logic [31:0] stage_6_out_10;
     logic [31:0] stage_6_out_11;
     logic [31:0] stage_6_out_12;
     logic [31:0] stage_6_out_13;
     logic [31:0] stage_6_out_14;
     logic [31:0] stage_6_out_15;
     logic [31:0] stage_6_out_16;
     logic [31:0] stage_6_out_17;
     logic [31:0] stage_6_out_18;
     logic [31:0] stage_6_out_19;
     logic [31:0] stage_6_out_20;
     logic [31:0] stage_6_out_21;
     logic [31:0] stage_6_out_22;
     logic [31:0] stage_6_out_23;
     logic [31:0] stage_6_out_24;
     logic [31:0] stage_6_out_25;
     logic [31:0] stage_6_out_26;
     logic [31:0] stage_6_out_27;
     logic [31:0] stage_6_out_28;
     logic [31:0] stage_6_out_29;
     logic [31:0] stage_6_out_30;
     logic [31:0] stage_6_out_31;
     logic [31:0] stage_6_out_32;
     logic [31:0] stage_6_out_33;
     logic [31:0] stage_7_out_0;
     logic [31:0] stage_7_out_1;
     logic [31:0] stage_7_out_2;
     logic [31:0] stage_7_out_3;
     logic [31:0] stage_7_out_4;
     logic [31:0] stage_7_out_5;
     logic [31:0] stage_7_out_6;
     logic [31:0] stage_7_out_7;
     logic [31:0] stage_7_out_8;
     logic [31:0] stage_7_out_9;
     logic [31:0] stage_7_out_10;
     logic [31:0] stage_7_out_11;
     logic [31:0] stage_7_out_12;
     logic [31:0] stage_7_out_13;
     logic [31:0] stage_7_out_14;
     logic [31:0] stage_7_out_15;
     logic [31:0] stage_7_out_16;
     logic [31:0] stage_7_out_17;
     logic [31:0] stage_7_out_18;
     logic [31:0] stage_7_out_19;
     logic [31:0] stage_7_out_20;
     logic [31:0] stage_7_out_21;
     logic [31:0] stage_7_out_22;
     logic [31:0] stage_7_out_23;
     logic [31:0] stage_7_out_24;
     logic [31:0] stage_7_out_25;
     logic [31:0] stage_7_out_26;
     logic [31:0] stage_7_out_27;
     logic [31:0] stage_7_out_28;
     logic [31:0] stage_7_out_29;
     logic [31:0] stage_7_out_30;
     logic [31:0] stage_7_out_31;
     logic [31:0] stage_7_out_32;
     logic [31:0] stage_7_out_33;
     logic [31:0] stage_8_out_0;
     logic [31:0] stage_8_out_1;
     logic [31:0] stage_8_out_2;
     logic [31:0] stage_8_out_3;
     logic [31:0] stage_8_out_4;
     logic [31:0] stage_8_out_5;
     logic [31:0] stage_8_out_6;
     logic [31:0] stage_8_out_7;
     logic [31:0] stage_8_out_8;
     logic [31:0] stage_8_out_9;
     logic [31:0] stage_8_out_10;
     logic [31:0] stage_8_out_11;
     logic [31:0] stage_8_out_12;
     logic [31:0] stage_8_out_13;
     logic [31:0] stage_8_out_14;
     logic [31:0] stage_8_out_15;
     logic [31:0] stage_8_out_16;
     logic [31:0] stage_8_out_17;
     logic [31:0] stage_8_out_18;
     logic [31:0] stage_8_out_19;
     logic [31:0] stage_8_out_20;
     logic [31:0] stage_8_out_21;
     logic [31:0] stage_8_out_22;
     logic [31:0] stage_8_out_23;
     logic [31:0] stage_8_out_24;
     logic [31:0] stage_8_out_25;
     logic [31:0] stage_8_out_26;
     logic [31:0] stage_8_out_27;
     logic [31:0] stage_8_out_28;
     logic [31:0] stage_8_out_29;
     logic [31:0] stage_8_out_30;
     logic [31:0] stage_8_out_31;
     logic [31:0] stage_8_out_32;
     logic [31:0] stage_8_out_33;
     logic [31:0] stage_9_out_0;
     logic [31:0] stage_9_out_1;
     logic [31:0] stage_9_out_2;
     logic [31:0] stage_9_out_3;
     logic [31:0] stage_9_out_4;
     logic [31:0] stage_9_out_5;
     logic [31:0] stage_9_out_6;
     logic [31:0] stage_9_out_7;
     logic [31:0] stage_9_out_8;
     logic [31:0] stage_9_out_9;
     logic [31:0] stage_9_out_10;
     logic [31:0] stage_9_out_11;
     logic [31:0] stage_9_out_12;
     logic [31:0] stage_9_out_13;
     logic [31:0] stage_9_out_14;
     logic [31:0] stage_9_out_15;
     logic [31:0] stage_9_out_16;
     logic [31:0] stage_9_out_17;
     logic [31:0] stage_9_out_18;
     logic [31:0] stage_9_out_19;
     logic [31:0] stage_9_out_20;
     logic [31:0] stage_9_out_21;
     logic [31:0] stage_9_out_22;
     logic [31:0] stage_9_out_23;
     logic [31:0] stage_9_out_24;
     logic [31:0] stage_9_out_25;
     logic [31:0] stage_9_out_26;
     logic [31:0] stage_9_out_27;
     logic [31:0] stage_9_out_28;
     logic [31:0] stage_9_out_29;
     logic [31:0] stage_9_out_30;
     logic [31:0] stage_9_out_31;
     logic [31:0] stage_9_out_32;
     logic [31:0] stage_9_out_33;
     logic [31:0] stage_10_out_0;
     logic [31:0] stage_10_out_1;
     logic [31:0] stage_10_out_2;
     logic [31:0] stage_10_out_3;
     logic [31:0] stage_10_out_4;
     logic [31:0] stage_10_out_5;
     logic [31:0] stage_10_out_6;
     logic [31:0] stage_10_out_7;
     logic [31:0] stage_10_out_8;
     logic [31:0] stage_10_out_9;
     logic [31:0] stage_10_out_10;
     logic [31:0] stage_10_out_11;
     logic [31:0] stage_10_out_12;
     logic [31:0] stage_10_out_13;
     logic [31:0] stage_10_out_14;
     logic [31:0] stage_10_out_15;
     logic [31:0] stage_10_out_16;
     logic [31:0] stage_10_out_17;
     logic [31:0] stage_10_out_18;
     logic [31:0] stage_10_out_19;
     logic [31:0] stage_10_out_20;
     logic [31:0] stage_10_out_21;
     logic [31:0] stage_10_out_22;
     logic [31:0] stage_10_out_23;
     logic [31:0] stage_10_out_24;
     logic [31:0] stage_10_out_25;
     logic [31:0] stage_10_out_26;
     logic [31:0] stage_10_out_27;
     logic [31:0] stage_10_out_28;
     logic [31:0] stage_10_out_29;
     logic [31:0] stage_10_out_30;
     logic [31:0] stage_10_out_31;
     logic [31:0] stage_10_out_32;
     logic [31:0] stage_10_out_33;
     logic [31:0] stage_11_out_0;
     logic [31:0] stage_11_out_1;
     logic [31:0] stage_11_out_2;
     logic [31:0] stage_11_out_3;
     logic [31:0] stage_11_out_4;
     logic [31:0] stage_11_out_5;
     logic [31:0] stage_11_out_6;
     logic [31:0] stage_11_out_7;
     logic [31:0] stage_11_out_8;
     logic [31:0] stage_11_out_9;
     logic [31:0] stage_11_out_10;
     logic [31:0] stage_11_out_11;
     logic [31:0] stage_11_out_12;
     logic [31:0] stage_11_out_13;
     logic [31:0] stage_11_out_14;
     logic [31:0] stage_11_out_15;
     logic [31:0] stage_11_out_16;
     logic [31:0] stage_11_out_17;
     logic [31:0] stage_11_out_18;
     logic [31:0] stage_11_out_19;
     logic [31:0] stage_11_out_20;
     logic [31:0] stage_11_out_21;
     logic [31:0] stage_11_out_22;
     logic [31:0] stage_11_out_23;
     logic [31:0] stage_11_out_24;
     logic [31:0] stage_11_out_25;
     logic [31:0] stage_11_out_26;
     logic [31:0] stage_11_out_27;
     logic [31:0] stage_11_out_28;
     logic [31:0] stage_11_out_29;
     logic [31:0] stage_11_out_30;
     logic [31:0] stage_11_out_31;
     logic [31:0] stage_11_out_32;
     logic [31:0] stage_11_out_33;
     logic [31:0] stage_12_out_0;
     logic [31:0] stage_12_out_1;
     logic [31:0] stage_12_out_2;
     logic [31:0] stage_12_out_3;
     logic [31:0] stage_12_out_4;
     logic [31:0] stage_12_out_5;
     logic [31:0] stage_12_out_6;
     logic [31:0] stage_12_out_7;
     logic [31:0] stage_12_out_8;
     logic [31:0] stage_12_out_9;
     logic [31:0] stage_12_out_10;
     logic [31:0] stage_12_out_11;
     logic [31:0] stage_12_out_12;
     logic [31:0] stage_12_out_13;
     logic [31:0] stage_12_out_14;
     logic [31:0] stage_12_out_15;
     logic [31:0] stage_12_out_16;
     logic [31:0] stage_12_out_17;
     logic [31:0] stage_12_out_18;
     logic [31:0] stage_12_out_19;
     logic [31:0] stage_12_out_20;
     logic [31:0] stage_12_out_21;
     logic [31:0] stage_12_out_22;
     logic [31:0] stage_12_out_23;
     logic [31:0] stage_12_out_24;
     logic [31:0] stage_12_out_25;
     logic [31:0] stage_12_out_26;
     logic [31:0] stage_12_out_27;
     logic [31:0] stage_12_out_28;
     logic [31:0] stage_12_out_29;
     logic [31:0] stage_12_out_30;
     logic [31:0] stage_12_out_31;
     logic [31:0] stage_12_out_32;
     logic [31:0] stage_12_out_33;
     logic [31:0] stage_13_out_0;
     logic [31:0] stage_13_out_1;
     logic [31:0] stage_13_out_2;
     logic [31:0] stage_13_out_3;
     logic [31:0] stage_13_out_4;
     logic [31:0] stage_13_out_5;
     logic [31:0] stage_13_out_6;
     logic [31:0] stage_13_out_7;
     logic [31:0] stage_13_out_8;
     logic [31:0] stage_13_out_9;
     logic [31:0] stage_13_out_10;
     logic [31:0] stage_13_out_11;
     logic [31:0] stage_13_out_12;
     logic [31:0] stage_13_out_13;
     logic [31:0] stage_13_out_14;
     logic [31:0] stage_13_out_15;
     logic [31:0] stage_13_out_16;
     logic [31:0] stage_13_out_17;
     logic [31:0] stage_13_out_18;
     logic [31:0] stage_13_out_19;
     logic [31:0] stage_13_out_20;
     logic [31:0] stage_13_out_21;
     logic [31:0] stage_13_out_22;
     logic [31:0] stage_13_out_23;
     logic [31:0] stage_13_out_24;
     logic [31:0] stage_13_out_25;
     logic [31:0] stage_13_out_26;
     logic [31:0] stage_13_out_27;
     logic [31:0] stage_13_out_28;
     logic [31:0] stage_13_out_29;
     logic [31:0] stage_13_out_30;
     logic [31:0] stage_13_out_31;
     logic [31:0] stage_13_out_32;
     logic [31:0] stage_13_out_33;
     logic [31:0] stage_14_out_0;
     logic [31:0] stage_14_out_1;
     logic [31:0] stage_14_out_2;
     logic [31:0] stage_14_out_3;
     logic [31:0] stage_14_out_4;
     logic [31:0] stage_14_out_5;
     logic [31:0] stage_14_out_6;
     logic [31:0] stage_14_out_7;
     logic [31:0] stage_14_out_8;
     logic [31:0] stage_14_out_9;
     logic [31:0] stage_14_out_10;
     logic [31:0] stage_14_out_11;
     logic [31:0] stage_14_out_12;
     logic [31:0] stage_14_out_13;
     logic [31:0] stage_14_out_14;
     logic [31:0] stage_14_out_15;
     logic [31:0] stage_14_out_16;
     logic [31:0] stage_14_out_17;
     logic [31:0] stage_14_out_18;
     logic [31:0] stage_14_out_19;
     logic [31:0] stage_14_out_20;
     logic [31:0] stage_14_out_21;
     logic [31:0] stage_14_out_22;
     logic [31:0] stage_14_out_23;
     logic [31:0] stage_14_out_24;
     logic [31:0] stage_14_out_25;
     logic [31:0] stage_14_out_26;
     logic [31:0] stage_14_out_27;
     logic [31:0] stage_14_out_28;
     logic [31:0] stage_14_out_29;
     logic [31:0] stage_14_out_30;
     logic [31:0] stage_14_out_31;
     logic [31:0] stage_14_out_32;
     logic [31:0] stage_14_out_33;
     logic [31:0] stage_15_out_0;
     logic [31:0] stage_15_out_1;
     logic [31:0] stage_15_out_2;
     logic [31:0] stage_15_out_3;
     logic [31:0] stage_15_out_4;
     logic [31:0] stage_15_out_5;
     logic [31:0] stage_15_out_6;
     logic [31:0] stage_15_out_7;
     logic [31:0] stage_15_out_8;
     logic [31:0] stage_15_out_9;
     logic [31:0] stage_15_out_10;
     logic [31:0] stage_15_out_11;
     logic [31:0] stage_15_out_12;
     logic [31:0] stage_15_out_13;
     logic [31:0] stage_15_out_14;
     logic [31:0] stage_15_out_15;
     logic [31:0] stage_15_out_16;
     logic [31:0] stage_15_out_17;
     logic [31:0] stage_15_out_18;
     logic [31:0] stage_15_out_19;
     logic [31:0] stage_15_out_20;
     logic [31:0] stage_15_out_21;
     logic [31:0] stage_15_out_22;
     logic [31:0] stage_15_out_23;
     logic [31:0] stage_15_out_24;
     logic [31:0] stage_15_out_25;
     logic [31:0] stage_15_out_26;
     logic [31:0] stage_15_out_27;
     logic [31:0] stage_15_out_28;
     logic [31:0] stage_15_out_29;
     logic [31:0] stage_15_out_30;
     logic [31:0] stage_15_out_31;
     logic [31:0] stage_15_out_32;
     logic [31:0] stage_15_out_33;
     logic [31:0] stage_16_out_0;
     logic [31:0] stage_16_out_1;
     logic [31:0] stage_16_out_2;
     logic [31:0] stage_16_out_3;
     logic [31:0] stage_16_out_4;
     logic [31:0] stage_16_out_5;
     logic [31:0] stage_16_out_6;
     logic [31:0] stage_16_out_7;
     logic [31:0] stage_16_out_8;
     logic [31:0] stage_16_out_9;
     logic [31:0] stage_16_out_10;
     logic [31:0] stage_16_out_11;
     logic [31:0] stage_16_out_12;
     logic [31:0] stage_16_out_13;
     logic [31:0] stage_16_out_14;
     logic [31:0] stage_16_out_15;
     logic [31:0] stage_16_out_16;
     logic [31:0] stage_16_out_17;
     logic [31:0] stage_16_out_18;
     logic [31:0] stage_16_out_19;
     logic [31:0] stage_16_out_20;
     logic [31:0] stage_16_out_21;
     logic [31:0] stage_16_out_22;
     logic [31:0] stage_16_out_23;
     logic [31:0] stage_16_out_24;
     logic [31:0] stage_16_out_25;
     logic [31:0] stage_16_out_26;
     logic [31:0] stage_16_out_27;
     logic [31:0] stage_16_out_28;
     logic [31:0] stage_16_out_29;
     logic [31:0] stage_16_out_30;
     logic [31:0] stage_16_out_31;
     logic [31:0] stage_16_out_32;
     logic [31:0] stage_16_out_33;
    assign stage_0_out_0 = (data_0 <= data_33) ? data_0 : data_33;
    assign stage_0_out_33 = (data_0 <= data_33) ? data_33 : data_0;
    assign stage_0_out_1 = (data_1 <= data_2) ? data_1 : data_2;
    assign stage_0_out_2 = (data_1 <= data_2) ? data_2 : data_1;
    assign stage_0_out_3 = (data_3 <= data_4) ? data_3 : data_4;
    assign stage_0_out_4 = (data_3 <= data_4) ? data_4 : data_3;
    assign stage_0_out_5 = (data_5 <= data_6) ? data_5 : data_6;
    assign stage_0_out_6 = (data_5 <= data_6) ? data_6 : data_5;
    assign stage_0_out_7 = (data_7 <= data_8) ? data_7 : data_8;
    assign stage_0_out_8 = (data_7 <= data_8) ? data_8 : data_7;
    assign stage_0_out_9 = (data_9 <= data_10) ? data_9 : data_10;
    assign stage_0_out_10 = (data_9 <= data_10) ? data_10 : data_9;
    assign stage_0_out_11 = (data_11 <= data_12) ? data_11 : data_12;
    assign stage_0_out_12 = (data_11 <= data_12) ? data_12 : data_11;
    assign stage_0_out_13 = (data_13 <= data_14) ? data_13 : data_14;
    assign stage_0_out_14 = (data_13 <= data_14) ? data_14 : data_13;
    assign stage_0_out_15 = (data_15 <= data_16) ? data_15 : data_16;
    assign stage_0_out_16 = (data_15 <= data_16) ? data_16 : data_15;
    assign stage_0_out_17 = (data_17 <= data_18) ? data_17 : data_18;
    assign stage_0_out_18 = (data_17 <= data_18) ? data_18 : data_17;
    assign stage_0_out_19 = (data_19 <= data_20) ? data_19 : data_20;
    assign stage_0_out_20 = (data_19 <= data_20) ? data_20 : data_19;
    assign stage_0_out_21 = (data_21 <= data_22) ? data_21 : data_22;
    assign stage_0_out_22 = (data_21 <= data_22) ? data_22 : data_21;
    assign stage_0_out_23 = (data_23 <= data_24) ? data_23 : data_24;
    assign stage_0_out_24 = (data_23 <= data_24) ? data_24 : data_23;
    assign stage_0_out_25 = (data_25 <= data_26) ? data_25 : data_26;
    assign stage_0_out_26 = (data_25 <= data_26) ? data_26 : data_25;
    assign stage_0_out_27 = (data_27 <= data_28) ? data_27 : data_28;
    assign stage_0_out_28 = (data_27 <= data_28) ? data_28 : data_27;
    assign stage_0_out_29 = (data_29 <= data_30) ? data_29 : data_30;
    assign stage_0_out_30 = (data_29 <= data_30) ? data_30 : data_29;
    assign stage_0_out_31 = (data_31 <= data_32) ? data_31 : data_32;
    assign stage_0_out_32 = (data_31 <= data_32) ? data_32 : data_31;
    assign stage_1_out_1 = (stage_0_out_1 <= stage_0_out_3) ? stage_0_out_1 : stage_0_out_3;
    assign stage_1_out_3 = (stage_0_out_1 <= stage_0_out_3) ? stage_0_out_3 : stage_0_out_1;
    assign stage_1_out_2 = (stage_0_out_2 <= stage_0_out_4) ? stage_0_out_2 : stage_0_out_4;
    assign stage_1_out_4 = (stage_0_out_2 <= stage_0_out_4) ? stage_0_out_4 : stage_0_out_2;
    assign stage_1_out_5 = (stage_0_out_5 <= stage_0_out_7) ? stage_0_out_5 : stage_0_out_7;
    assign stage_1_out_7 = (stage_0_out_5 <= stage_0_out_7) ? stage_0_out_7 : stage_0_out_5;
    assign stage_1_out_6 = (stage_0_out_6 <= stage_0_out_8) ? stage_0_out_6 : stage_0_out_8;
    assign stage_1_out_8 = (stage_0_out_6 <= stage_0_out_8) ? stage_0_out_8 : stage_0_out_6;
    assign stage_1_out_9 = (stage_0_out_9 <= stage_0_out_11) ? stage_0_out_9 : stage_0_out_11;
    assign stage_1_out_11 = (stage_0_out_9 <= stage_0_out_11) ? stage_0_out_11 : stage_0_out_9;
    assign stage_1_out_10 = (stage_0_out_10 <= stage_0_out_12) ? stage_0_out_10 : stage_0_out_12;
    assign stage_1_out_12 = (stage_0_out_10 <= stage_0_out_12) ? stage_0_out_12 : stage_0_out_10;
    assign stage_1_out_13 = (stage_0_out_13 <= stage_0_out_15) ? stage_0_out_13 : stage_0_out_15;
    assign stage_1_out_15 = (stage_0_out_13 <= stage_0_out_15) ? stage_0_out_15 : stage_0_out_13;
    assign stage_1_out_14 = (stage_0_out_14 <= stage_0_out_16) ? stage_0_out_14 : stage_0_out_16;
    assign stage_1_out_16 = (stage_0_out_14 <= stage_0_out_16) ? stage_0_out_16 : stage_0_out_14;
    assign stage_1_out_17 = (stage_0_out_17 <= stage_0_out_19) ? stage_0_out_17 : stage_0_out_19;
    assign stage_1_out_19 = (stage_0_out_17 <= stage_0_out_19) ? stage_0_out_19 : stage_0_out_17;
    assign stage_1_out_18 = (stage_0_out_18 <= stage_0_out_20) ? stage_0_out_18 : stage_0_out_20;
    assign stage_1_out_20 = (stage_0_out_18 <= stage_0_out_20) ? stage_0_out_20 : stage_0_out_18;
    assign stage_1_out_21 = (stage_0_out_21 <= stage_0_out_23) ? stage_0_out_21 : stage_0_out_23;
    assign stage_1_out_23 = (stage_0_out_21 <= stage_0_out_23) ? stage_0_out_23 : stage_0_out_21;
    assign stage_1_out_22 = (stage_0_out_22 <= stage_0_out_24) ? stage_0_out_22 : stage_0_out_24;
    assign stage_1_out_24 = (stage_0_out_22 <= stage_0_out_24) ? stage_0_out_24 : stage_0_out_22;
    assign stage_1_out_25 = (stage_0_out_25 <= stage_0_out_27) ? stage_0_out_25 : stage_0_out_27;
    assign stage_1_out_27 = (stage_0_out_25 <= stage_0_out_27) ? stage_0_out_27 : stage_0_out_25;
    assign stage_1_out_26 = (stage_0_out_26 <= stage_0_out_28) ? stage_0_out_26 : stage_0_out_28;
    assign stage_1_out_28 = (stage_0_out_26 <= stage_0_out_28) ? stage_0_out_28 : stage_0_out_26;
    assign stage_1_out_29 = (stage_0_out_29 <= stage_0_out_31) ? stage_0_out_29 : stage_0_out_31;
    assign stage_1_out_31 = (stage_0_out_29 <= stage_0_out_31) ? stage_0_out_31 : stage_0_out_29;
    assign stage_1_out_30 = (stage_0_out_30 <= stage_0_out_32) ? stage_0_out_30 : stage_0_out_32;
    assign stage_1_out_32 = (stage_0_out_30 <= stage_0_out_32) ? stage_0_out_32 : stage_0_out_30;
    assign stage_1_out_0 = stage_0_out_0;
    assign stage_1_out_33 = stage_0_out_33;
    assign stage_2_out_1 = (stage_1_out_1 <= stage_1_out_5) ? stage_1_out_1 : stage_1_out_5;
    assign stage_2_out_5 = (stage_1_out_1 <= stage_1_out_5) ? stage_1_out_5 : stage_1_out_1;
    assign stage_2_out_2 = (stage_1_out_2 <= stage_1_out_6) ? stage_1_out_2 : stage_1_out_6;
    assign stage_2_out_6 = (stage_1_out_2 <= stage_1_out_6) ? stage_1_out_6 : stage_1_out_2;
    assign stage_2_out_3 = (stage_1_out_3 <= stage_1_out_7) ? stage_1_out_3 : stage_1_out_7;
    assign stage_2_out_7 = (stage_1_out_3 <= stage_1_out_7) ? stage_1_out_7 : stage_1_out_3;
    assign stage_2_out_4 = (stage_1_out_4 <= stage_1_out_8) ? stage_1_out_4 : stage_1_out_8;
    assign stage_2_out_8 = (stage_1_out_4 <= stage_1_out_8) ? stage_1_out_8 : stage_1_out_4;
    assign stage_2_out_9 = (stage_1_out_9 <= stage_1_out_13) ? stage_1_out_9 : stage_1_out_13;
    assign stage_2_out_13 = (stage_1_out_9 <= stage_1_out_13) ? stage_1_out_13 : stage_1_out_9;
    assign stage_2_out_10 = (stage_1_out_10 <= stage_1_out_14) ? stage_1_out_10 : stage_1_out_14;
    assign stage_2_out_14 = (stage_1_out_10 <= stage_1_out_14) ? stage_1_out_14 : stage_1_out_10;
    assign stage_2_out_11 = (stage_1_out_11 <= stage_1_out_15) ? stage_1_out_11 : stage_1_out_15;
    assign stage_2_out_15 = (stage_1_out_11 <= stage_1_out_15) ? stage_1_out_15 : stage_1_out_11;
    assign stage_2_out_12 = (stage_1_out_12 <= stage_1_out_16) ? stage_1_out_12 : stage_1_out_16;
    assign stage_2_out_16 = (stage_1_out_12 <= stage_1_out_16) ? stage_1_out_16 : stage_1_out_12;
    assign stage_2_out_17 = (stage_1_out_17 <= stage_1_out_21) ? stage_1_out_17 : stage_1_out_21;
    assign stage_2_out_21 = (stage_1_out_17 <= stage_1_out_21) ? stage_1_out_21 : stage_1_out_17;
    assign stage_2_out_18 = (stage_1_out_18 <= stage_1_out_22) ? stage_1_out_18 : stage_1_out_22;
    assign stage_2_out_22 = (stage_1_out_18 <= stage_1_out_22) ? stage_1_out_22 : stage_1_out_18;
    assign stage_2_out_19 = (stage_1_out_19 <= stage_1_out_23) ? stage_1_out_19 : stage_1_out_23;
    assign stage_2_out_23 = (stage_1_out_19 <= stage_1_out_23) ? stage_1_out_23 : stage_1_out_19;
    assign stage_2_out_20 = (stage_1_out_20 <= stage_1_out_24) ? stage_1_out_20 : stage_1_out_24;
    assign stage_2_out_24 = (stage_1_out_20 <= stage_1_out_24) ? stage_1_out_24 : stage_1_out_20;
    assign stage_2_out_25 = (stage_1_out_25 <= stage_1_out_29) ? stage_1_out_25 : stage_1_out_29;
    assign stage_2_out_29 = (stage_1_out_25 <= stage_1_out_29) ? stage_1_out_29 : stage_1_out_25;
    assign stage_2_out_26 = (stage_1_out_26 <= stage_1_out_30) ? stage_1_out_26 : stage_1_out_30;
    assign stage_2_out_30 = (stage_1_out_26 <= stage_1_out_30) ? stage_1_out_30 : stage_1_out_26;
    assign stage_2_out_27 = (stage_1_out_27 <= stage_1_out_31) ? stage_1_out_27 : stage_1_out_31;
    assign stage_2_out_31 = (stage_1_out_27 <= stage_1_out_31) ? stage_1_out_31 : stage_1_out_27;
    assign stage_2_out_28 = (stage_1_out_28 <= stage_1_out_32) ? stage_1_out_28 : stage_1_out_32;
    assign stage_2_out_32 = (stage_1_out_28 <= stage_1_out_32) ? stage_1_out_32 : stage_1_out_28;
    assign stage_2_out_0 = stage_1_out_0;
    assign stage_2_out_33 = stage_1_out_33;
    assign stage_3_out_1 = (stage_2_out_1 <= stage_2_out_9) ? stage_2_out_1 : stage_2_out_9;
    assign stage_3_out_9 = (stage_2_out_1 <= stage_2_out_9) ? stage_2_out_9 : stage_2_out_1;
    assign stage_3_out_2 = (stage_2_out_2 <= stage_2_out_10) ? stage_2_out_2 : stage_2_out_10;
    assign stage_3_out_10 = (stage_2_out_2 <= stage_2_out_10) ? stage_2_out_10 : stage_2_out_2;
    assign stage_3_out_3 = (stage_2_out_3 <= stage_2_out_11) ? stage_2_out_3 : stage_2_out_11;
    assign stage_3_out_11 = (stage_2_out_3 <= stage_2_out_11) ? stage_2_out_11 : stage_2_out_3;
    assign stage_3_out_4 = (stage_2_out_4 <= stage_2_out_12) ? stage_2_out_4 : stage_2_out_12;
    assign stage_3_out_12 = (stage_2_out_4 <= stage_2_out_12) ? stage_2_out_12 : stage_2_out_4;
    assign stage_3_out_5 = (stage_2_out_5 <= stage_2_out_13) ? stage_2_out_5 : stage_2_out_13;
    assign stage_3_out_13 = (stage_2_out_5 <= stage_2_out_13) ? stage_2_out_13 : stage_2_out_5;
    assign stage_3_out_6 = (stage_2_out_6 <= stage_2_out_14) ? stage_2_out_6 : stage_2_out_14;
    assign stage_3_out_14 = (stage_2_out_6 <= stage_2_out_14) ? stage_2_out_14 : stage_2_out_6;
    assign stage_3_out_7 = (stage_2_out_7 <= stage_2_out_15) ? stage_2_out_7 : stage_2_out_15;
    assign stage_3_out_15 = (stage_2_out_7 <= stage_2_out_15) ? stage_2_out_15 : stage_2_out_7;
    assign stage_3_out_8 = (stage_2_out_8 <= stage_2_out_16) ? stage_2_out_8 : stage_2_out_16;
    assign stage_3_out_16 = (stage_2_out_8 <= stage_2_out_16) ? stage_2_out_16 : stage_2_out_8;
    assign stage_3_out_17 = (stage_2_out_17 <= stage_2_out_25) ? stage_2_out_17 : stage_2_out_25;
    assign stage_3_out_25 = (stage_2_out_17 <= stage_2_out_25) ? stage_2_out_25 : stage_2_out_17;
    assign stage_3_out_18 = (stage_2_out_18 <= stage_2_out_26) ? stage_2_out_18 : stage_2_out_26;
    assign stage_3_out_26 = (stage_2_out_18 <= stage_2_out_26) ? stage_2_out_26 : stage_2_out_18;
    assign stage_3_out_19 = (stage_2_out_19 <= stage_2_out_27) ? stage_2_out_19 : stage_2_out_27;
    assign stage_3_out_27 = (stage_2_out_19 <= stage_2_out_27) ? stage_2_out_27 : stage_2_out_19;
    assign stage_3_out_20 = (stage_2_out_20 <= stage_2_out_28) ? stage_2_out_20 : stage_2_out_28;
    assign stage_3_out_28 = (stage_2_out_20 <= stage_2_out_28) ? stage_2_out_28 : stage_2_out_20;
    assign stage_3_out_21 = (stage_2_out_21 <= stage_2_out_29) ? stage_2_out_21 : stage_2_out_29;
    assign stage_3_out_29 = (stage_2_out_21 <= stage_2_out_29) ? stage_2_out_29 : stage_2_out_21;
    assign stage_3_out_22 = (stage_2_out_22 <= stage_2_out_30) ? stage_2_out_22 : stage_2_out_30;
    assign stage_3_out_30 = (stage_2_out_22 <= stage_2_out_30) ? stage_2_out_30 : stage_2_out_22;
    assign stage_3_out_23 = (stage_2_out_23 <= stage_2_out_31) ? stage_2_out_23 : stage_2_out_31;
    assign stage_3_out_31 = (stage_2_out_23 <= stage_2_out_31) ? stage_2_out_31 : stage_2_out_23;
    assign stage_3_out_24 = (stage_2_out_24 <= stage_2_out_32) ? stage_2_out_24 : stage_2_out_32;
    assign stage_3_out_32 = (stage_2_out_24 <= stage_2_out_32) ? stage_2_out_32 : stage_2_out_24;
    assign stage_3_out_0 = stage_2_out_0;
    assign stage_3_out_33 = stage_2_out_33;
    assign stage_4_out_1 = (stage_3_out_1 <= stage_3_out_17) ? stage_3_out_1 : stage_3_out_17;
    assign stage_4_out_17 = (stage_3_out_1 <= stage_3_out_17) ? stage_3_out_17 : stage_3_out_1;
    assign stage_4_out_2 = (stage_3_out_2 <= stage_3_out_18) ? stage_3_out_2 : stage_3_out_18;
    assign stage_4_out_18 = (stage_3_out_2 <= stage_3_out_18) ? stage_3_out_18 : stage_3_out_2;
    assign stage_4_out_3 = (stage_3_out_3 <= stage_3_out_19) ? stage_3_out_3 : stage_3_out_19;
    assign stage_4_out_19 = (stage_3_out_3 <= stage_3_out_19) ? stage_3_out_19 : stage_3_out_3;
    assign stage_4_out_4 = (stage_3_out_4 <= stage_3_out_20) ? stage_3_out_4 : stage_3_out_20;
    assign stage_4_out_20 = (stage_3_out_4 <= stage_3_out_20) ? stage_3_out_20 : stage_3_out_4;
    assign stage_4_out_5 = (stage_3_out_5 <= stage_3_out_21) ? stage_3_out_5 : stage_3_out_21;
    assign stage_4_out_21 = (stage_3_out_5 <= stage_3_out_21) ? stage_3_out_21 : stage_3_out_5;
    assign stage_4_out_6 = (stage_3_out_6 <= stage_3_out_22) ? stage_3_out_6 : stage_3_out_22;
    assign stage_4_out_22 = (stage_3_out_6 <= stage_3_out_22) ? stage_3_out_22 : stage_3_out_6;
    assign stage_4_out_7 = (stage_3_out_7 <= stage_3_out_23) ? stage_3_out_7 : stage_3_out_23;
    assign stage_4_out_23 = (stage_3_out_7 <= stage_3_out_23) ? stage_3_out_23 : stage_3_out_7;
    assign stage_4_out_8 = (stage_3_out_8 <= stage_3_out_24) ? stage_3_out_8 : stage_3_out_24;
    assign stage_4_out_24 = (stage_3_out_8 <= stage_3_out_24) ? stage_3_out_24 : stage_3_out_8;
    assign stage_4_out_9 = (stage_3_out_9 <= stage_3_out_25) ? stage_3_out_9 : stage_3_out_25;
    assign stage_4_out_25 = (stage_3_out_9 <= stage_3_out_25) ? stage_3_out_25 : stage_3_out_9;
    assign stage_4_out_10 = (stage_3_out_10 <= stage_3_out_26) ? stage_3_out_10 : stage_3_out_26;
    assign stage_4_out_26 = (stage_3_out_10 <= stage_3_out_26) ? stage_3_out_26 : stage_3_out_10;
    assign stage_4_out_11 = (stage_3_out_11 <= stage_3_out_27) ? stage_3_out_11 : stage_3_out_27;
    assign stage_4_out_27 = (stage_3_out_11 <= stage_3_out_27) ? stage_3_out_27 : stage_3_out_11;
    assign stage_4_out_12 = (stage_3_out_12 <= stage_3_out_28) ? stage_3_out_12 : stage_3_out_28;
    assign stage_4_out_28 = (stage_3_out_12 <= stage_3_out_28) ? stage_3_out_28 : stage_3_out_12;
    assign stage_4_out_13 = (stage_3_out_13 <= stage_3_out_29) ? stage_3_out_13 : stage_3_out_29;
    assign stage_4_out_29 = (stage_3_out_13 <= stage_3_out_29) ? stage_3_out_29 : stage_3_out_13;
    assign stage_4_out_14 = (stage_3_out_14 <= stage_3_out_30) ? stage_3_out_14 : stage_3_out_30;
    assign stage_4_out_30 = (stage_3_out_14 <= stage_3_out_30) ? stage_3_out_30 : stage_3_out_14;
    assign stage_4_out_15 = (stage_3_out_15 <= stage_3_out_31) ? stage_3_out_15 : stage_3_out_31;
    assign stage_4_out_31 = (stage_3_out_15 <= stage_3_out_31) ? stage_3_out_31 : stage_3_out_15;
    assign stage_4_out_16 = (stage_3_out_16 <= stage_3_out_32) ? stage_3_out_16 : stage_3_out_32;
    assign stage_4_out_32 = (stage_3_out_16 <= stage_3_out_32) ? stage_3_out_32 : stage_3_out_16;
    assign stage_4_out_0 = stage_3_out_0;
    assign stage_4_out_33 = stage_3_out_33;
    assign stage_5_out_0 = (stage_4_out_0 <= stage_4_out_4) ? stage_4_out_0 : stage_4_out_4;
    assign stage_5_out_4 = (stage_4_out_0 <= stage_4_out_4) ? stage_4_out_4 : stage_4_out_0;
    assign stage_5_out_2 = (stage_4_out_2 <= stage_4_out_3) ? stage_4_out_2 : stage_4_out_3;
    assign stage_5_out_3 = (stage_4_out_2 <= stage_4_out_3) ? stage_4_out_3 : stage_4_out_2;
    assign stage_5_out_5 = (stage_4_out_5 <= stage_4_out_17) ? stage_4_out_5 : stage_4_out_17;
    assign stage_5_out_17 = (stage_4_out_5 <= stage_4_out_17) ? stage_4_out_17 : stage_4_out_5;
    assign stage_5_out_6 = (stage_4_out_6 <= stage_4_out_11) ? stage_4_out_6 : stage_4_out_11;
    assign stage_5_out_11 = (stage_4_out_6 <= stage_4_out_11) ? stage_4_out_11 : stage_4_out_6;
    assign stage_5_out_7 = (stage_4_out_7 <= stage_4_out_10) ? stage_4_out_7 : stage_4_out_10;
    assign stage_5_out_10 = (stage_4_out_7 <= stage_4_out_10) ? stage_4_out_10 : stage_4_out_7;
    assign stage_5_out_8 = (stage_4_out_8 <= stage_4_out_12) ? stage_4_out_8 : stage_4_out_12;
    assign stage_5_out_12 = (stage_4_out_8 <= stage_4_out_12) ? stage_4_out_12 : stage_4_out_8;
    assign stage_5_out_14 = (stage_4_out_14 <= stage_4_out_15) ? stage_4_out_14 : stage_4_out_15;
    assign stage_5_out_15 = (stage_4_out_14 <= stage_4_out_15) ? stage_4_out_15 : stage_4_out_14;
    assign stage_5_out_16 = (stage_4_out_16 <= stage_4_out_28) ? stage_4_out_16 : stage_4_out_28;
    assign stage_5_out_28 = (stage_4_out_16 <= stage_4_out_28) ? stage_4_out_28 : stage_4_out_16;
    assign stage_5_out_18 = (stage_4_out_18 <= stage_4_out_19) ? stage_4_out_18 : stage_4_out_19;
    assign stage_5_out_19 = (stage_4_out_18 <= stage_4_out_19) ? stage_4_out_19 : stage_4_out_18;
    assign stage_5_out_21 = (stage_4_out_21 <= stage_4_out_25) ? stage_4_out_21 : stage_4_out_25;
    assign stage_5_out_25 = (stage_4_out_21 <= stage_4_out_25) ? stage_4_out_25 : stage_4_out_21;
    assign stage_5_out_22 = (stage_4_out_22 <= stage_4_out_27) ? stage_4_out_22 : stage_4_out_27;
    assign stage_5_out_27 = (stage_4_out_22 <= stage_4_out_27) ? stage_4_out_27 : stage_4_out_22;
    assign stage_5_out_23 = (stage_4_out_23 <= stage_4_out_26) ? stage_4_out_23 : stage_4_out_26;
    assign stage_5_out_26 = (stage_4_out_23 <= stage_4_out_26) ? stage_4_out_26 : stage_4_out_23;
    assign stage_5_out_29 = (stage_4_out_29 <= stage_4_out_33) ? stage_4_out_29 : stage_4_out_33;
    assign stage_5_out_33 = (stage_4_out_29 <= stage_4_out_33) ? stage_4_out_33 : stage_4_out_29;
    assign stage_5_out_30 = (stage_4_out_30 <= stage_4_out_31) ? stage_4_out_30 : stage_4_out_31;
    assign stage_5_out_31 = (stage_4_out_30 <= stage_4_out_31) ? stage_4_out_31 : stage_4_out_30;
    assign stage_5_out_1 = stage_4_out_1;
    assign stage_5_out_9 = stage_4_out_9;
    assign stage_5_out_13 = stage_4_out_13;
    assign stage_5_out_20 = stage_4_out_20;
    assign stage_5_out_24 = stage_4_out_24;
    assign stage_5_out_32 = stage_4_out_32;
    assign stage_6_out_0 = (stage_5_out_0 <= stage_5_out_7) ? stage_5_out_0 : stage_5_out_7;
    assign stage_6_out_7 = (stage_5_out_0 <= stage_5_out_7) ? stage_5_out_7 : stage_5_out_0;
    assign stage_6_out_2 = (stage_5_out_2 <= stage_5_out_9) ? stage_5_out_2 : stage_5_out_9;
    assign stage_6_out_9 = (stage_5_out_2 <= stage_5_out_9) ? stage_5_out_9 : stage_5_out_2;
    assign stage_6_out_4 = (stage_5_out_4 <= stage_5_out_13) ? stage_5_out_4 : stage_5_out_13;
    assign stage_6_out_13 = (stage_5_out_4 <= stage_5_out_13) ? stage_5_out_13 : stage_5_out_4;
    assign stage_6_out_8 = (stage_5_out_8 <= stage_5_out_14) ? stage_5_out_8 : stage_5_out_14;
    assign stage_6_out_14 = (stage_5_out_8 <= stage_5_out_14) ? stage_5_out_14 : stage_5_out_8;
    assign stage_6_out_19 = (stage_5_out_19 <= stage_5_out_25) ? stage_5_out_19 : stage_5_out_25;
    assign stage_6_out_25 = (stage_5_out_19 <= stage_5_out_25) ? stage_5_out_25 : stage_5_out_19;
    assign stage_6_out_20 = (stage_5_out_20 <= stage_5_out_29) ? stage_5_out_20 : stage_5_out_29;
    assign stage_6_out_29 = (stage_5_out_20 <= stage_5_out_29) ? stage_5_out_29 : stage_5_out_20;
    assign stage_6_out_24 = (stage_5_out_24 <= stage_5_out_31) ? stage_5_out_24 : stage_5_out_31;
    assign stage_6_out_31 = (stage_5_out_24 <= stage_5_out_31) ? stage_5_out_31 : stage_5_out_24;
    assign stage_6_out_26 = (stage_5_out_26 <= stage_5_out_33) ? stage_5_out_26 : stage_5_out_33;
    assign stage_6_out_33 = (stage_5_out_26 <= stage_5_out_33) ? stage_5_out_33 : stage_5_out_26;
    assign stage_6_out_6 = (stage_5_out_6 <= stage_5_out_10) ? stage_5_out_6 : stage_5_out_10;
    assign stage_6_out_10 = (stage_5_out_6 <= stage_5_out_10) ? stage_5_out_10 : stage_5_out_6;
    assign stage_6_out_12 = (stage_5_out_12 <= stage_5_out_15) ? stage_5_out_12 : stage_5_out_15;
    assign stage_6_out_15 = (stage_5_out_12 <= stage_5_out_15) ? stage_5_out_15 : stage_5_out_12;
    assign stage_6_out_18 = (stage_5_out_18 <= stage_5_out_21) ? stage_5_out_18 : stage_5_out_21;
    assign stage_6_out_21 = (stage_5_out_18 <= stage_5_out_21) ? stage_5_out_21 : stage_5_out_18;
    assign stage_6_out_23 = (stage_5_out_23 <= stage_5_out_27) ? stage_5_out_23 : stage_5_out_27;
    assign stage_6_out_27 = (stage_5_out_23 <= stage_5_out_27) ? stage_5_out_27 : stage_5_out_23;
    assign stage_6_out_3 = (stage_5_out_3 <= stage_5_out_5) ? stage_5_out_3 : stage_5_out_5;
    assign stage_6_out_5 = (stage_5_out_3 <= stage_5_out_5) ? stage_5_out_5 : stage_5_out_3;
    assign stage_6_out_28 = (stage_5_out_28 <= stage_5_out_30) ? stage_5_out_28 : stage_5_out_30;
    assign stage_6_out_30 = (stage_5_out_28 <= stage_5_out_30) ? stage_5_out_30 : stage_5_out_28;
    assign stage_6_out_11 = (stage_5_out_11 <= stage_5_out_17) ? stage_5_out_11 : stage_5_out_17;
    assign stage_6_out_17 = (stage_5_out_11 <= stage_5_out_17) ? stage_5_out_17 : stage_5_out_11;
    assign stage_6_out_16 = (stage_5_out_16 <= stage_5_out_22) ? stage_5_out_16 : stage_5_out_22;
    assign stage_6_out_22 = (stage_5_out_16 <= stage_5_out_22) ? stage_5_out_22 : stage_5_out_16;
    assign stage_6_out_1 = stage_5_out_1;
    assign stage_6_out_32 = stage_5_out_32;
    assign stage_7_out_0 = (stage_6_out_0 <= stage_6_out_9) ? stage_6_out_0 : stage_6_out_9;
    assign stage_7_out_9 = (stage_6_out_0 <= stage_6_out_9) ? stage_6_out_9 : stage_6_out_0;
    assign stage_7_out_4 = (stage_6_out_4 <= stage_6_out_18) ? stage_6_out_4 : stage_6_out_18;
    assign stage_7_out_18 = (stage_6_out_4 <= stage_6_out_18) ? stage_6_out_18 : stage_6_out_4;
    assign stage_7_out_7 = (stage_6_out_7 <= stage_6_out_21) ? stage_6_out_7 : stage_6_out_21;
    assign stage_7_out_21 = (stage_6_out_7 <= stage_6_out_21) ? stage_6_out_21 : stage_6_out_7;
    assign stage_7_out_8 = (stage_6_out_8 <= stage_6_out_19) ? stage_6_out_8 : stage_6_out_19;
    assign stage_7_out_19 = (stage_6_out_8 <= stage_6_out_19) ? stage_6_out_19 : stage_6_out_8;
    assign stage_7_out_10 = (stage_6_out_10 <= stage_6_out_20) ? stage_6_out_10 : stage_6_out_20;
    assign stage_7_out_20 = (stage_6_out_10 <= stage_6_out_20) ? stage_6_out_20 : stage_6_out_10;
    assign stage_7_out_12 = (stage_6_out_12 <= stage_6_out_26) ? stage_6_out_12 : stage_6_out_26;
    assign stage_7_out_26 = (stage_6_out_12 <= stage_6_out_26) ? stage_6_out_26 : stage_6_out_12;
    assign stage_7_out_13 = (stage_6_out_13 <= stage_6_out_23) ? stage_6_out_13 : stage_6_out_23;
    assign stage_7_out_23 = (stage_6_out_13 <= stage_6_out_23) ? stage_6_out_23 : stage_6_out_13;
    assign stage_7_out_14 = (stage_6_out_14 <= stage_6_out_25) ? stage_6_out_14 : stage_6_out_25;
    assign stage_7_out_25 = (stage_6_out_14 <= stage_6_out_25) ? stage_6_out_25 : stage_6_out_14;
    assign stage_7_out_15 = (stage_6_out_15 <= stage_6_out_29) ? stage_6_out_15 : stage_6_out_29;
    assign stage_7_out_29 = (stage_6_out_15 <= stage_6_out_29) ? stage_6_out_29 : stage_6_out_15;
    assign stage_7_out_24 = (stage_6_out_24 <= stage_6_out_33) ? stage_6_out_24 : stage_6_out_33;
    assign stage_7_out_33 = (stage_6_out_24 <= stage_6_out_33) ? stage_6_out_33 : stage_6_out_24;
    assign stage_7_out_16 = (stage_6_out_16 <= stage_6_out_17) ? stage_6_out_16 : stage_6_out_17;
    assign stage_7_out_17 = (stage_6_out_16 <= stage_6_out_17) ? stage_6_out_17 : stage_6_out_16;
    assign stage_7_out_1 = stage_6_out_1;
    assign stage_7_out_2 = stage_6_out_2;
    assign stage_7_out_3 = stage_6_out_3;
    assign stage_7_out_5 = stage_6_out_5;
    assign stage_7_out_6 = stage_6_out_6;
    assign stage_7_out_11 = stage_6_out_11;
    assign stage_7_out_22 = stage_6_out_22;
    assign stage_7_out_27 = stage_6_out_27;
    assign stage_7_out_28 = stage_6_out_28;
    assign stage_7_out_30 = stage_6_out_30;
    assign stage_7_out_31 = stage_6_out_31;
    assign stage_7_out_32 = stage_6_out_32;
    assign stage_8_out_33 = (stage_7_out_33 <= stage_7_out_28) ? stage_7_out_33 : stage_7_out_28;
    assign stage_8_out_28 = (stage_7_out_33 <= stage_7_out_28) ? stage_7_out_28 : stage_7_out_33;
    assign stage_8_out_24 = (stage_7_out_24 <= stage_7_out_16) ? stage_7_out_24 : stage_7_out_16;
    assign stage_8_out_16 = (stage_7_out_24 <= stage_7_out_16) ? stage_7_out_16 : stage_7_out_24;
    assign stage_8_out_22 = (stage_7_out_22 <= stage_7_out_13) ? stage_7_out_22 : stage_7_out_13;
    assign stage_8_out_13 = (stage_7_out_22 <= stage_7_out_13) ? stage_7_out_13 : stage_7_out_22;
    assign stage_8_out_20 = (stage_7_out_20 <= stage_7_out_11) ? stage_7_out_20 : stage_7_out_11;
    assign stage_8_out_11 = (stage_7_out_20 <= stage_7_out_11) ? stage_7_out_11 : stage_7_out_20;
    assign stage_8_out_17 = (stage_7_out_17 <= stage_7_out_9) ? stage_7_out_17 : stage_7_out_9;
    assign stage_8_out_9 = (stage_7_out_17 <= stage_7_out_9) ? stage_7_out_9 : stage_7_out_17;
    assign stage_8_out_5 = (stage_7_out_5 <= stage_7_out_0) ? stage_7_out_5 : stage_7_out_0;
    assign stage_8_out_0 = (stage_7_out_5 <= stage_7_out_0) ? stage_7_out_0 : stage_7_out_5;
    assign stage_8_out_29 = (stage_7_out_29 <= stage_7_out_27) ? stage_7_out_29 : stage_7_out_27;
    assign stage_8_out_27 = (stage_7_out_29 <= stage_7_out_27) ? stage_7_out_27 : stage_7_out_29;
    assign stage_8_out_6 = (stage_7_out_6 <= stage_7_out_4) ? stage_7_out_6 : stage_7_out_4;
    assign stage_8_out_4 = (stage_7_out_6 <= stage_7_out_4) ? stage_7_out_4 : stage_7_out_6;
    assign stage_8_out_25 = (stage_7_out_25 <= stage_7_out_23) ? stage_7_out_25 : stage_7_out_23;
    assign stage_8_out_23 = (stage_7_out_25 <= stage_7_out_23) ? stage_7_out_23 : stage_7_out_25;
    assign stage_8_out_10 = (stage_7_out_10 <= stage_7_out_8) ? stage_7_out_10 : stage_7_out_8;
    assign stage_8_out_8 = (stage_7_out_10 <= stage_7_out_8) ? stage_7_out_8 : stage_7_out_10;
    assign stage_8_out_21 = (stage_7_out_21 <= stage_7_out_15) ? stage_7_out_21 : stage_7_out_15;
    assign stage_8_out_15 = (stage_7_out_21 <= stage_7_out_15) ? stage_7_out_15 : stage_7_out_21;
    assign stage_8_out_18 = (stage_7_out_18 <= stage_7_out_12) ? stage_7_out_18 : stage_7_out_12;
    assign stage_8_out_12 = (stage_7_out_18 <= stage_7_out_12) ? stage_7_out_12 : stage_7_out_18;
    assign stage_9_out_33 = (stage_8_out_33 <= stage_8_out_24) ? stage_8_out_33 : stage_8_out_24;
    assign stage_9_out_24 = (stage_8_out_33 <= stage_8_out_24) ? stage_8_out_24 : stage_8_out_33;
    assign stage_9_out_29 = (stage_8_out_29 <= stage_8_out_15) ? stage_8_out_29 : stage_8_out_15;
    assign stage_9_out_15 = (stage_8_out_29 <= stage_8_out_15) ? stage_8_out_15 : stage_8_out_29;
    assign stage_9_out_26 = (stage_8_out_26 <= stage_8_out_12) ? stage_8_out_26 : stage_8_out_12;
    assign stage_9_out_12 = (stage_8_out_26 <= stage_8_out_12) ? stage_8_out_12 : stage_8_out_26;
    assign stage_9_out_25 = (stage_8_out_25 <= stage_8_out_14) ? stage_8_out_25 : stage_8_out_14;
    assign stage_9_out_14 = (stage_8_out_25 <= stage_8_out_14) ? stage_8_out_14 : stage_8_out_25;
    assign stage_9_out_23 = (stage_8_out_23 <= stage_8_out_13) ? stage_8_out_23 : stage_8_out_13;
    assign stage_9_out_13 = (stage_8_out_23 <= stage_8_out_13) ? stage_8_out_13 : stage_8_out_23;
    assign stage_9_out_21 = (stage_8_out_21 <= stage_8_out_7) ? stage_8_out_21 : stage_8_out_7;
    assign stage_9_out_7 = (stage_8_out_21 <= stage_8_out_7) ? stage_8_out_7 : stage_8_out_21;
    assign stage_9_out_20 = (stage_8_out_20 <= stage_8_out_10) ? stage_8_out_20 : stage_8_out_10;
    assign stage_9_out_10 = (stage_8_out_20 <= stage_8_out_10) ? stage_8_out_10 : stage_8_out_20;
    assign stage_9_out_19 = (stage_8_out_19 <= stage_8_out_8) ? stage_8_out_19 : stage_8_out_8;
    assign stage_9_out_8 = (stage_8_out_19 <= stage_8_out_8) ? stage_8_out_8 : stage_8_out_19;
    assign stage_9_out_18 = (stage_8_out_18 <= stage_8_out_4) ? stage_8_out_18 : stage_8_out_4;
    assign stage_9_out_4 = (stage_8_out_18 <= stage_8_out_4) ? stage_8_out_4 : stage_8_out_18;
    assign stage_9_out_9 = (stage_8_out_9 <= stage_8_out_0) ? stage_8_out_9 : stage_8_out_0;
    assign stage_9_out_0 = (stage_8_out_9 <= stage_8_out_0) ? stage_8_out_0 : stage_8_out_9;
    assign stage_9_out_17 = (stage_8_out_17 <= stage_8_out_16) ? stage_8_out_17 : stage_8_out_16;
    assign stage_9_out_16 = (stage_8_out_17 <= stage_8_out_16) ? stage_8_out_16 : stage_8_out_17;
    assign stage_10_out_33 = (stage_9_out_33 <= stage_9_out_26) ? stage_9_out_33 : stage_9_out_26;
    assign stage_10_out_26 = (stage_9_out_33 <= stage_9_out_26) ? stage_9_out_26 : stage_9_out_33;
    assign stage_10_out_31 = (stage_9_out_31 <= stage_9_out_24) ? stage_9_out_31 : stage_9_out_24;
    assign stage_10_out_24 = (stage_9_out_31 <= stage_9_out_24) ? stage_9_out_24 : stage_9_out_31;
    assign stage_10_out_29 = (stage_9_out_29 <= stage_9_out_20) ? stage_9_out_29 : stage_9_out_20;
    assign stage_10_out_20 = (stage_9_out_29 <= stage_9_out_20) ? stage_9_out_20 : stage_9_out_29;
    assign stage_10_out_25 = (stage_9_out_25 <= stage_9_out_19) ? stage_9_out_25 : stage_9_out_19;
    assign stage_10_out_19 = (stage_9_out_25 <= stage_9_out_19) ? stage_9_out_19 : stage_9_out_25;
    assign stage_10_out_14 = (stage_9_out_14 <= stage_9_out_8) ? stage_9_out_14 : stage_9_out_8;
    assign stage_10_out_8 = (stage_9_out_14 <= stage_9_out_8) ? stage_9_out_8 : stage_9_out_14;
    assign stage_10_out_13 = (stage_9_out_13 <= stage_9_out_4) ? stage_9_out_13 : stage_9_out_4;
    assign stage_10_out_4 = (stage_9_out_13 <= stage_9_out_4) ? stage_9_out_4 : stage_9_out_13;
    assign stage_10_out_9 = (stage_9_out_9 <= stage_9_out_2) ? stage_9_out_9 : stage_9_out_2;
    assign stage_10_out_2 = (stage_9_out_9 <= stage_9_out_2) ? stage_9_out_2 : stage_9_out_9;
    assign stage_10_out_7 = (stage_9_out_7 <= stage_9_out_0) ? stage_9_out_7 : stage_9_out_0;
    assign stage_10_out_0 = (stage_9_out_7 <= stage_9_out_0) ? stage_9_out_0 : stage_9_out_7;
    assign stage_10_out_27 = (stage_9_out_27 <= stage_9_out_23) ? stage_9_out_27 : stage_9_out_23;
    assign stage_10_out_23 = (stage_9_out_27 <= stage_9_out_23) ? stage_9_out_23 : stage_9_out_27;
    assign stage_10_out_21 = (stage_9_out_21 <= stage_9_out_18) ? stage_9_out_21 : stage_9_out_18;
    assign stage_10_out_18 = (stage_9_out_21 <= stage_9_out_18) ? stage_9_out_18 : stage_9_out_21;
    assign stage_10_out_15 = (stage_9_out_15 <= stage_9_out_12) ? stage_9_out_15 : stage_9_out_12;
    assign stage_10_out_12 = (stage_9_out_15 <= stage_9_out_12) ? stage_9_out_12 : stage_9_out_15;
    assign stage_10_out_10 = (stage_9_out_10 <= stage_9_out_6) ? stage_9_out_10 : stage_9_out_6;
    assign stage_10_out_6 = (stage_9_out_10 <= stage_9_out_6) ? stage_9_out_6 : stage_9_out_10;
    assign stage_10_out_30 = (stage_9_out_30 <= stage_9_out_28) ? stage_9_out_30 : stage_9_out_28;
    assign stage_10_out_28 = (stage_9_out_30 <= stage_9_out_28) ? stage_9_out_28 : stage_9_out_30;
    assign stage_10_out_5 = (stage_9_out_5 <= stage_9_out_3) ? stage_9_out_5 : stage_9_out_3;
    assign stage_10_out_3 = (stage_9_out_5 <= stage_9_out_3) ? stage_9_out_3 : stage_9_out_5;
    assign stage_10_out_22 = (stage_9_out_22 <= stage_9_out_16) ? stage_9_out_22 : stage_9_out_16;
    assign stage_10_out_16 = (stage_9_out_22 <= stage_9_out_16) ? stage_9_out_16 : stage_9_out_22;
    assign stage_10_out_17 = (stage_9_out_17 <= stage_9_out_11) ? stage_9_out_17 : stage_9_out_11;
    assign stage_10_out_11 = (stage_9_out_17 <= stage_9_out_11) ? stage_9_out_11 : stage_9_out_17;
    assign stage_11_out_33 = (stage_10_out_33 <= stage_10_out_29) ? stage_10_out_33 : stage_10_out_29;
    assign stage_11_out_29 = (stage_10_out_33 <= stage_10_out_29) ? stage_10_out_29 : stage_10_out_33;
    assign stage_11_out_31 = (stage_10_out_31 <= stage_10_out_30) ? stage_10_out_31 : stage_10_out_30;
    assign stage_11_out_30 = (stage_10_out_31 <= stage_10_out_30) ? stage_10_out_30 : stage_10_out_31;
    assign stage_11_out_28 = (stage_10_out_28 <= stage_10_out_16) ? stage_10_out_28 : stage_10_out_16;
    assign stage_11_out_16 = (stage_10_out_28 <= stage_10_out_16) ? stage_10_out_16 : stage_10_out_28;
    assign stage_11_out_27 = (stage_10_out_27 <= stage_10_out_22) ? stage_10_out_27 : stage_10_out_22;
    assign stage_11_out_22 = (stage_10_out_27 <= stage_10_out_22) ? stage_10_out_22 : stage_10_out_27;
    assign stage_11_out_26 = (stage_10_out_26 <= stage_10_out_23) ? stage_10_out_26 : stage_10_out_23;
    assign stage_11_out_23 = (stage_10_out_26 <= stage_10_out_23) ? stage_10_out_23 : stage_10_out_26;
    assign stage_11_out_25 = (stage_10_out_25 <= stage_10_out_21) ? stage_10_out_25 : stage_10_out_21;
    assign stage_11_out_21 = (stage_10_out_25 <= stage_10_out_21) ? stage_10_out_21 : stage_10_out_25;
    assign stage_11_out_19 = (stage_10_out_19 <= stage_10_out_18) ? stage_10_out_19 : stage_10_out_18;
    assign stage_11_out_18 = (stage_10_out_19 <= stage_10_out_18) ? stage_10_out_18 : stage_10_out_19;
    assign stage_11_out_17 = (stage_10_out_17 <= stage_10_out_5) ? stage_10_out_17 : stage_10_out_5;
    assign stage_11_out_5 = (stage_10_out_17 <= stage_10_out_5) ? stage_10_out_5 : stage_10_out_17;
    assign stage_11_out_15 = (stage_10_out_15 <= stage_10_out_14) ? stage_10_out_15 : stage_10_out_14;
    assign stage_11_out_14 = (stage_10_out_15 <= stage_10_out_14) ? stage_10_out_14 : stage_10_out_15;
    assign stage_11_out_12 = (stage_10_out_12 <= stage_10_out_8) ? stage_10_out_12 : stage_10_out_8;
    assign stage_11_out_8 = (stage_10_out_12 <= stage_10_out_8) ? stage_10_out_8 : stage_10_out_12;
    assign stage_11_out_11 = (stage_10_out_11 <= stage_10_out_6) ? stage_10_out_11 : stage_10_out_6;
    assign stage_11_out_6 = (stage_10_out_11 <= stage_10_out_6) ? stage_10_out_6 : stage_10_out_11;
    assign stage_11_out_10 = (stage_10_out_10 <= stage_10_out_7) ? stage_10_out_10 : stage_10_out_7;
    assign stage_11_out_7 = (stage_10_out_10 <= stage_10_out_7) ? stage_10_out_7 : stage_10_out_10;
    assign stage_11_out_4 = (stage_10_out_4 <= stage_10_out_0) ? stage_10_out_4 : stage_10_out_0;
    assign stage_11_out_0 = (stage_10_out_4 <= stage_10_out_0) ? stage_10_out_0 : stage_10_out_4;
    assign stage_11_out_3 = (stage_10_out_3 <= stage_10_out_2) ? stage_10_out_3 : stage_10_out_2;
    assign stage_11_out_2 = (stage_10_out_3 <= stage_10_out_2) ? stage_10_out_2 : stage_10_out_3;
    assign stage_12_out_32 = (stage_11_out_32 <= stage_11_out_16) ? stage_11_out_32 : stage_11_out_16;
    assign stage_12_out_16 = (stage_11_out_32 <= stage_11_out_16) ? stage_11_out_16 : stage_11_out_32;
    assign stage_12_out_31 = (stage_11_out_31 <= stage_11_out_15) ? stage_11_out_31 : stage_11_out_15;
    assign stage_12_out_15 = (stage_11_out_31 <= stage_11_out_15) ? stage_11_out_15 : stage_11_out_31;
    assign stage_12_out_30 = (stage_11_out_30 <= stage_11_out_14) ? stage_11_out_30 : stage_11_out_14;
    assign stage_12_out_14 = (stage_11_out_30 <= stage_11_out_14) ? stage_11_out_14 : stage_11_out_30;
    assign stage_12_out_29 = (stage_11_out_29 <= stage_11_out_13) ? stage_11_out_29 : stage_11_out_13;
    assign stage_12_out_13 = (stage_11_out_29 <= stage_11_out_13) ? stage_11_out_13 : stage_11_out_29;
    assign stage_12_out_28 = (stage_11_out_28 <= stage_11_out_12) ? stage_11_out_28 : stage_11_out_12;
    assign stage_12_out_12 = (stage_11_out_28 <= stage_11_out_12) ? stage_11_out_12 : stage_11_out_28;
    assign stage_12_out_27 = (stage_11_out_27 <= stage_11_out_11) ? stage_11_out_27 : stage_11_out_11;
    assign stage_12_out_11 = (stage_11_out_27 <= stage_11_out_11) ? stage_11_out_11 : stage_11_out_27;
    assign stage_12_out_26 = (stage_11_out_26 <= stage_11_out_10) ? stage_11_out_26 : stage_11_out_10;
    assign stage_12_out_10 = (stage_11_out_26 <= stage_11_out_10) ? stage_11_out_10 : stage_11_out_26;
    assign stage_12_out_25 = (stage_11_out_25 <= stage_11_out_9) ? stage_11_out_25 : stage_11_out_9;
    assign stage_12_out_9 = (stage_11_out_25 <= stage_11_out_9) ? stage_11_out_9 : stage_11_out_25;
    assign stage_12_out_24 = (stage_11_out_24 <= stage_11_out_8) ? stage_11_out_24 : stage_11_out_8;
    assign stage_12_out_8 = (stage_11_out_24 <= stage_11_out_8) ? stage_11_out_8 : stage_11_out_24;
    assign stage_12_out_23 = (stage_11_out_23 <= stage_11_out_7) ? stage_11_out_23 : stage_11_out_7;
    assign stage_12_out_7 = (stage_11_out_23 <= stage_11_out_7) ? stage_11_out_7 : stage_11_out_23;
    assign stage_12_out_22 = (stage_11_out_22 <= stage_11_out_6) ? stage_11_out_22 : stage_11_out_6;
    assign stage_12_out_6 = (stage_11_out_22 <= stage_11_out_6) ? stage_11_out_6 : stage_11_out_22;
    assign stage_12_out_21 = (stage_11_out_21 <= stage_11_out_5) ? stage_11_out_21 : stage_11_out_5;
    assign stage_12_out_5 = (stage_11_out_21 <= stage_11_out_5) ? stage_11_out_5 : stage_11_out_21;
    assign stage_12_out_20 = (stage_11_out_20 <= stage_11_out_4) ? stage_11_out_20 : stage_11_out_4;
    assign stage_12_out_4 = (stage_11_out_20 <= stage_11_out_4) ? stage_11_out_4 : stage_11_out_20;
    assign stage_12_out_19 = (stage_11_out_19 <= stage_11_out_3) ? stage_11_out_19 : stage_11_out_3;
    assign stage_12_out_3 = (stage_11_out_19 <= stage_11_out_3) ? stage_11_out_3 : stage_11_out_19;
    assign stage_12_out_18 = (stage_11_out_18 <= stage_11_out_2) ? stage_11_out_18 : stage_11_out_2;
    assign stage_12_out_2 = (stage_11_out_18 <= stage_11_out_2) ? stage_11_out_2 : stage_11_out_18;
    assign stage_12_out_17 = (stage_11_out_17 <= stage_11_out_1) ? stage_11_out_17 : stage_11_out_1;
    assign stage_12_out_1 = (stage_11_out_17 <= stage_11_out_1) ? stage_11_out_1 : stage_11_out_17;
    assign stage_13_out_32 = (stage_12_out_32 <= stage_12_out_24) ? stage_12_out_32 : stage_12_out_24;
    assign stage_13_out_24 = (stage_12_out_32 <= stage_12_out_24) ? stage_12_out_24 : stage_12_out_32;
    assign stage_13_out_31 = (stage_12_out_31 <= stage_12_out_23) ? stage_12_out_31 : stage_12_out_23;
    assign stage_13_out_23 = (stage_12_out_31 <= stage_12_out_23) ? stage_12_out_23 : stage_12_out_31;
    assign stage_13_out_30 = (stage_12_out_30 <= stage_12_out_22) ? stage_12_out_30 : stage_12_out_22;
    assign stage_13_out_22 = (stage_12_out_30 <= stage_12_out_22) ? stage_12_out_22 : stage_12_out_30;
    assign stage_13_out_29 = (stage_12_out_29 <= stage_12_out_21) ? stage_12_out_29 : stage_12_out_21;
    assign stage_13_out_21 = (stage_12_out_29 <= stage_12_out_21) ? stage_12_out_21 : stage_12_out_29;
    assign stage_13_out_28 = (stage_12_out_28 <= stage_12_out_20) ? stage_12_out_28 : stage_12_out_20;
    assign stage_13_out_20 = (stage_12_out_28 <= stage_12_out_20) ? stage_12_out_20 : stage_12_out_28;
    assign stage_13_out_27 = (stage_12_out_27 <= stage_12_out_19) ? stage_12_out_27 : stage_12_out_19;
    assign stage_13_out_19 = (stage_12_out_27 <= stage_12_out_19) ? stage_12_out_19 : stage_12_out_27;
    assign stage_13_out_26 = (stage_12_out_26 <= stage_12_out_18) ? stage_12_out_26 : stage_12_out_18;
    assign stage_13_out_18 = (stage_12_out_26 <= stage_12_out_18) ? stage_12_out_18 : stage_12_out_26;
    assign stage_13_out_25 = (stage_12_out_25 <= stage_12_out_17) ? stage_12_out_25 : stage_12_out_17;
    assign stage_13_out_17 = (stage_12_out_25 <= stage_12_out_17) ? stage_12_out_17 : stage_12_out_25;
    assign stage_13_out_16 = (stage_12_out_16 <= stage_12_out_8) ? stage_12_out_16 : stage_12_out_8;
    assign stage_13_out_8 = (stage_12_out_16 <= stage_12_out_8) ? stage_12_out_8 : stage_12_out_16;
    assign stage_13_out_15 = (stage_12_out_15 <= stage_12_out_7) ? stage_12_out_15 : stage_12_out_7;
    assign stage_13_out_7 = (stage_12_out_15 <= stage_12_out_7) ? stage_12_out_7 : stage_12_out_15;
    assign stage_13_out_14 = (stage_12_out_14 <= stage_12_out_6) ? stage_12_out_14 : stage_12_out_6;
    assign stage_13_out_6 = (stage_12_out_14 <= stage_12_out_6) ? stage_12_out_6 : stage_12_out_14;
    assign stage_13_out_13 = (stage_12_out_13 <= stage_12_out_5) ? stage_12_out_13 : stage_12_out_5;
    assign stage_13_out_5 = (stage_12_out_13 <= stage_12_out_5) ? stage_12_out_5 : stage_12_out_13;
    assign stage_13_out_12 = (stage_12_out_12 <= stage_12_out_4) ? stage_12_out_12 : stage_12_out_4;
    assign stage_13_out_4 = (stage_12_out_12 <= stage_12_out_4) ? stage_12_out_4 : stage_12_out_12;
    assign stage_13_out_11 = (stage_12_out_11 <= stage_12_out_3) ? stage_12_out_11 : stage_12_out_3;
    assign stage_13_out_3 = (stage_12_out_11 <= stage_12_out_3) ? stage_12_out_3 : stage_12_out_11;
    assign stage_13_out_10 = (stage_12_out_10 <= stage_12_out_2) ? stage_12_out_10 : stage_12_out_2;
    assign stage_13_out_2 = (stage_12_out_10 <= stage_12_out_2) ? stage_12_out_2 : stage_12_out_10;
    assign stage_13_out_9 = (stage_12_out_9 <= stage_12_out_1) ? stage_12_out_9 : stage_12_out_1;
    assign stage_13_out_1 = (stage_12_out_9 <= stage_12_out_1) ? stage_12_out_1 : stage_12_out_9;
    assign stage_14_out_32 = (stage_13_out_32 <= stage_13_out_28) ? stage_13_out_32 : stage_13_out_28;
    assign stage_14_out_28 = (stage_13_out_32 <= stage_13_out_28) ? stage_13_out_28 : stage_13_out_32;
    assign stage_14_out_31 = (stage_13_out_31 <= stage_13_out_27) ? stage_13_out_31 : stage_13_out_27;
    assign stage_14_out_27 = (stage_13_out_31 <= stage_13_out_27) ? stage_13_out_27 : stage_13_out_31;
    assign stage_14_out_30 = (stage_13_out_30 <= stage_13_out_26) ? stage_13_out_30 : stage_13_out_26;
    assign stage_14_out_26 = (stage_13_out_30 <= stage_13_out_26) ? stage_13_out_26 : stage_13_out_30;
    assign stage_14_out_29 = (stage_13_out_29 <= stage_13_out_25) ? stage_13_out_29 : stage_13_out_25;
    assign stage_14_out_25 = (stage_13_out_29 <= stage_13_out_25) ? stage_13_out_25 : stage_13_out_29;
    assign stage_14_out_24 = (stage_13_out_24 <= stage_13_out_20) ? stage_13_out_24 : stage_13_out_20;
    assign stage_14_out_20 = (stage_13_out_24 <= stage_13_out_20) ? stage_13_out_20 : stage_13_out_24;
    assign stage_14_out_23 = (stage_13_out_23 <= stage_13_out_19) ? stage_13_out_23 : stage_13_out_19;
    assign stage_14_out_19 = (stage_13_out_23 <= stage_13_out_19) ? stage_13_out_19 : stage_13_out_23;
    assign stage_14_out_22 = (stage_13_out_22 <= stage_13_out_18) ? stage_13_out_22 : stage_13_out_18;
    assign stage_14_out_18 = (stage_13_out_22 <= stage_13_out_18) ? stage_13_out_18 : stage_13_out_22;
    assign stage_14_out_21 = (stage_13_out_21 <= stage_13_out_17) ? stage_13_out_21 : stage_13_out_17;
    assign stage_14_out_17 = (stage_13_out_21 <= stage_13_out_17) ? stage_13_out_17 : stage_13_out_21;
    assign stage_14_out_16 = (stage_13_out_16 <= stage_13_out_12) ? stage_13_out_16 : stage_13_out_12;
    assign stage_14_out_12 = (stage_13_out_16 <= stage_13_out_12) ? stage_13_out_12 : stage_13_out_16;
    assign stage_14_out_15 = (stage_13_out_15 <= stage_13_out_11) ? stage_13_out_15 : stage_13_out_11;
    assign stage_14_out_11 = (stage_13_out_15 <= stage_13_out_11) ? stage_13_out_11 : stage_13_out_15;
    assign stage_14_out_14 = (stage_13_out_14 <= stage_13_out_10) ? stage_13_out_14 : stage_13_out_10;
    assign stage_14_out_10 = (stage_13_out_14 <= stage_13_out_10) ? stage_13_out_10 : stage_13_out_14;
    assign stage_14_out_13 = (stage_13_out_13 <= stage_13_out_9) ? stage_13_out_13 : stage_13_out_9;
    assign stage_14_out_9 = (stage_13_out_13 <= stage_13_out_9) ? stage_13_out_9 : stage_13_out_13;
    assign stage_14_out_8 = (stage_13_out_8 <= stage_13_out_4) ? stage_13_out_8 : stage_13_out_4;
    assign stage_14_out_4 = (stage_13_out_8 <= stage_13_out_4) ? stage_13_out_4 : stage_13_out_8;
    assign stage_14_out_7 = (stage_13_out_7 <= stage_13_out_3) ? stage_13_out_7 : stage_13_out_3;
    assign stage_14_out_3 = (stage_13_out_7 <= stage_13_out_3) ? stage_13_out_3 : stage_13_out_7;
    assign stage_14_out_6 = (stage_13_out_6 <= stage_13_out_2) ? stage_13_out_6 : stage_13_out_2;
    assign stage_14_out_2 = (stage_13_out_6 <= stage_13_out_2) ? stage_13_out_2 : stage_13_out_6;
    assign stage_14_out_5 = (stage_13_out_5 <= stage_13_out_1) ? stage_13_out_5 : stage_13_out_1;
    assign stage_14_out_1 = (stage_13_out_5 <= stage_13_out_1) ? stage_13_out_1 : stage_13_out_5;
    assign stage_15_out_32 = (stage_14_out_32 <= stage_14_out_30) ? stage_14_out_32 : stage_14_out_30;
    assign stage_15_out_30 = (stage_14_out_32 <= stage_14_out_30) ? stage_14_out_30 : stage_14_out_32;
    assign stage_15_out_31 = (stage_14_out_31 <= stage_14_out_29) ? stage_14_out_31 : stage_14_out_29;
    assign stage_15_out_29 = (stage_14_out_31 <= stage_14_out_29) ? stage_14_out_29 : stage_14_out_31;
    assign stage_15_out_28 = (stage_14_out_28 <= stage_14_out_26) ? stage_14_out_28 : stage_14_out_26;
    assign stage_15_out_26 = (stage_14_out_28 <= stage_14_out_26) ? stage_14_out_26 : stage_14_out_28;
    assign stage_15_out_27 = (stage_14_out_27 <= stage_14_out_25) ? stage_14_out_27 : stage_14_out_25;
    assign stage_15_out_25 = (stage_14_out_27 <= stage_14_out_25) ? stage_14_out_25 : stage_14_out_27;
    assign stage_15_out_24 = (stage_14_out_24 <= stage_14_out_22) ? stage_14_out_24 : stage_14_out_22;
    assign stage_15_out_22 = (stage_14_out_24 <= stage_14_out_22) ? stage_14_out_22 : stage_14_out_24;
    assign stage_15_out_23 = (stage_14_out_23 <= stage_14_out_21) ? stage_14_out_23 : stage_14_out_21;
    assign stage_15_out_21 = (stage_14_out_23 <= stage_14_out_21) ? stage_14_out_21 : stage_14_out_23;
    assign stage_15_out_20 = (stage_14_out_20 <= stage_14_out_18) ? stage_14_out_20 : stage_14_out_18;
    assign stage_15_out_18 = (stage_14_out_20 <= stage_14_out_18) ? stage_14_out_18 : stage_14_out_20;
    assign stage_15_out_19 = (stage_14_out_19 <= stage_14_out_17) ? stage_14_out_19 : stage_14_out_17;
    assign stage_15_out_17 = (stage_14_out_19 <= stage_14_out_17) ? stage_14_out_17 : stage_14_out_19;
    assign stage_15_out_16 = (stage_14_out_16 <= stage_14_out_14) ? stage_14_out_16 : stage_14_out_14;
    assign stage_15_out_14 = (stage_14_out_16 <= stage_14_out_14) ? stage_14_out_14 : stage_14_out_16;
    assign stage_15_out_15 = (stage_14_out_15 <= stage_14_out_13) ? stage_14_out_15 : stage_14_out_13;
    assign stage_15_out_13 = (stage_14_out_15 <= stage_14_out_13) ? stage_14_out_13 : stage_14_out_15;
    assign stage_15_out_12 = (stage_14_out_12 <= stage_14_out_10) ? stage_14_out_12 : stage_14_out_10;
    assign stage_15_out_10 = (stage_14_out_12 <= stage_14_out_10) ? stage_14_out_10 : stage_14_out_12;
    assign stage_15_out_11 = (stage_14_out_11 <= stage_14_out_9) ? stage_14_out_11 : stage_14_out_9;
    assign stage_15_out_9 = (stage_14_out_11 <= stage_14_out_9) ? stage_14_out_9 : stage_14_out_11;
    assign stage_15_out_8 = (stage_14_out_8 <= stage_14_out_6) ? stage_14_out_8 : stage_14_out_6;
    assign stage_15_out_6 = (stage_14_out_8 <= stage_14_out_6) ? stage_14_out_6 : stage_14_out_8;
    assign stage_15_out_7 = (stage_14_out_7 <= stage_14_out_5) ? stage_14_out_7 : stage_14_out_5;
    assign stage_15_out_5 = (stage_14_out_7 <= stage_14_out_5) ? stage_14_out_5 : stage_14_out_7;
    assign stage_15_out_4 = (stage_14_out_4 <= stage_14_out_2) ? stage_14_out_4 : stage_14_out_2;
    assign stage_15_out_2 = (stage_14_out_4 <= stage_14_out_2) ? stage_14_out_2 : stage_14_out_4;
    assign stage_15_out_3 = (stage_14_out_3 <= stage_14_out_1) ? stage_14_out_3 : stage_14_out_1;
    assign stage_15_out_1 = (stage_14_out_3 <= stage_14_out_1) ? stage_14_out_1 : stage_14_out_3;
    assign stage_16_out_33 = (stage_15_out_33 <= stage_15_out_0) ? stage_15_out_33 : stage_15_out_0;
    assign stage_16_out_0 = (stage_15_out_33 <= stage_15_out_0) ? stage_15_out_0 : stage_15_out_33;
    assign stage_16_out_32 = (stage_15_out_32 <= stage_15_out_31) ? stage_15_out_32 : stage_15_out_31;
    assign stage_16_out_31 = (stage_15_out_32 <= stage_15_out_31) ? stage_15_out_31 : stage_15_out_32;
    assign stage_16_out_30 = (stage_15_out_30 <= stage_15_out_29) ? stage_15_out_30 : stage_15_out_29;
    assign stage_16_out_29 = (stage_15_out_30 <= stage_15_out_29) ? stage_15_out_29 : stage_15_out_30;
    assign stage_16_out_28 = (stage_15_out_28 <= stage_15_out_27) ? stage_15_out_28 : stage_15_out_27;
    assign stage_16_out_27 = (stage_15_out_28 <= stage_15_out_27) ? stage_15_out_27 : stage_15_out_28;
    assign stage_16_out_26 = (stage_15_out_26 <= stage_15_out_25) ? stage_15_out_26 : stage_15_out_25;
    assign stage_16_out_25 = (stage_15_out_26 <= stage_15_out_25) ? stage_15_out_25 : stage_15_out_26;
    assign stage_16_out_24 = (stage_15_out_24 <= stage_15_out_23) ? stage_15_out_24 : stage_15_out_23;
    assign stage_16_out_23 = (stage_15_out_24 <= stage_15_out_23) ? stage_15_out_23 : stage_15_out_24;
    assign stage_16_out_22 = (stage_15_out_22 <= stage_15_out_21) ? stage_15_out_22 : stage_15_out_21;
    assign stage_16_out_21 = (stage_15_out_22 <= stage_15_out_21) ? stage_15_out_21 : stage_15_out_22;
    assign stage_16_out_20 = (stage_15_out_20 <= stage_15_out_19) ? stage_15_out_20 : stage_15_out_19;
    assign stage_16_out_19 = (stage_15_out_20 <= stage_15_out_19) ? stage_15_out_19 : stage_15_out_20;
    assign stage_16_out_18 = (stage_15_out_18 <= stage_15_out_17) ? stage_15_out_18 : stage_15_out_17;
    assign stage_16_out_17 = (stage_15_out_18 <= stage_15_out_17) ? stage_15_out_17 : stage_15_out_18;
    assign stage_16_out_16 = (stage_15_out_16 <= stage_15_out_15) ? stage_15_out_16 : stage_15_out_15;
    assign stage_16_out_15 = (stage_15_out_16 <= stage_15_out_15) ? stage_15_out_15 : stage_15_out_16;
    assign stage_16_out_14 = (stage_15_out_14 <= stage_15_out_13) ? stage_15_out_14 : stage_15_out_13;
    assign stage_16_out_13 = (stage_15_out_14 <= stage_15_out_13) ? stage_15_out_13 : stage_15_out_14;
    assign stage_16_out_12 = (stage_15_out_12 <= stage_15_out_11) ? stage_15_out_12 : stage_15_out_11;
    assign stage_16_out_11 = (stage_15_out_12 <= stage_15_out_11) ? stage_15_out_11 : stage_15_out_12;
    assign stage_16_out_10 = (stage_15_out_10 <= stage_15_out_9) ? stage_15_out_10 : stage_15_out_9;
    assign stage_16_out_9 = (stage_15_out_10 <= stage_15_out_9) ? stage_15_out_9 : stage_15_out_10;
    assign stage_16_out_8 = (stage_15_out_8 <= stage_15_out_7) ? stage_15_out_8 : stage_15_out_7;
    assign stage_16_out_7 = (stage_15_out_8 <= stage_15_out_7) ? stage_15_out_7 : stage_15_out_8;
    assign stage_16_out_6 = (stage_15_out_6 <= stage_15_out_5) ? stage_15_out_6 : stage_15_out_5;
    assign stage_16_out_5 = (stage_15_out_6 <= stage_15_out_5) ? stage_15_out_5 : stage_15_out_6;
    assign stage_16_out_4 = (stage_15_out_4 <= stage_15_out_3) ? stage_15_out_4 : stage_15_out_3;
    assign stage_16_out_3 = (stage_15_out_4 <= stage_15_out_3) ? stage_15_out_3 : stage_15_out_4;
    assign stage_16_out_2 = (stage_15_out_2 <= stage_15_out_1) ? stage_15_out_2 : stage_15_out_1;
    assign stage_16_out_1 = (stage_15_out_2 <= stage_15_out_1) ? stage_15_out_1 : stage_15_out_2;
    assign sort_0 = stage_16_out_0;
    assign sort_1 = stage_16_out_1;
    assign sort_2 = stage_16_out_2;
    assign sort_3 = stage_16_out_3;
    assign sort_4 = stage_16_out_4;
    assign sort_5 = stage_16_out_5;
    assign sort_6 = stage_16_out_6;
    assign sort_7 = stage_16_out_7;
    assign sort_8 = stage_16_out_8;
    assign sort_9 = stage_16_out_9;
    assign sort_10 = stage_16_out_10;
    assign sort_11 = stage_16_out_11;
    assign sort_12 = stage_16_out_12;
    assign sort_13 = stage_16_out_13;
    assign sort_14 = stage_16_out_14;
    assign sort_15 = stage_16_out_15;
    assign sort_16 = stage_16_out_16;
    assign sort_17 = stage_16_out_17;
    assign sort_18 = stage_16_out_18;
    assign sort_19 = stage_16_out_19;
    assign sort_20 = stage_16_out_20;
    assign sort_21 = stage_16_out_21;
    assign sort_22 = stage_16_out_22;
    assign sort_23 = stage_16_out_23;
    assign sort_24 = stage_16_out_24;
    assign sort_25 = stage_16_out_25;
    assign sort_26 = stage_16_out_26;
    assign sort_27 = stage_16_out_27;
    assign sort_28 = stage_16_out_28;
    assign sort_29 = stage_16_out_29;
    assign sort_30 = stage_16_out_30;
    assign sort_31 = stage_16_out_31;
    assign sort_32 = stage_16_out_32;
    assign sort_33 = stage_16_out_33;
endmodule

module sort_34_209_17_tb;

    logic clk;
    data_t data_0;
    data_t data_1;
    data_t data_2;
    data_t data_3;
    data_t data_4;
    data_t data_5;
    data_t data_6;
    data_t data_7;
    data_t data_8;
    data_t data_9;
    data_t data_10;
    data_t data_11;
    data_t data_12;
    data_t data_13;
    data_t data_14;
    data_t data_15;
    data_t data_16;
    data_t data_17;
    data_t data_18;
    data_t data_19;
    data_t data_20;
    data_t data_21;
    data_t data_22;
    data_t data_23;
    data_t data_24;
    data_t data_25;
    data_t data_26;
    data_t data_27;
    data_t data_28;
    data_t data_29;
    data_t data_30;
    data_t data_31;
    data_t data_32;
    data_t data_33;
    data_t sort_0;
    data_t sort_1;
    data_t sort_2;
    data_t sort_3;
    data_t sort_4;
    data_t sort_5;
    data_t sort_6;
    data_t sort_7;
    data_t sort_8;
    data_t sort_9;
    data_t sort_10;
    data_t sort_11;
    data_t sort_12;
    data_t sort_13;
    data_t sort_14;
    data_t sort_15;
    data_t sort_16;
    data_t sort_17;
    data_t sort_18;
    data_t sort_19;
    data_t sort_20;
    data_t sort_21;
    data_t sort_22;
    data_t sort_23;
    data_t sort_24;
    data_t sort_25;
    data_t sort_26;
    data_t sort_27;
    data_t sort_28;
    data_t sort_29;
    data_t sort_30;
    data_t sort_31;
    data_t sort_32;
    data_t sort_33;

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Instantiate DUT
    sort_34_209_17 dut (
        .clk(clk),
        .data_0(data_0),
        .data_1(data_1),
        .data_2(data_2),
        .data_3(data_3),
        .data_4(data_4),
        .data_5(data_5),
        .data_6(data_6),
        .data_7(data_7),
        .data_8(data_8),
        .data_9(data_9),
        .data_10(data_10),
        .data_11(data_11),
        .data_12(data_12),
        .data_13(data_13),
        .data_14(data_14),
        .data_15(data_15),
        .data_16(data_16),
        .data_17(data_17),
        .data_18(data_18),
        .data_19(data_19),
        .data_20(data_20),
        .data_21(data_21),
        .data_22(data_22),
        .data_23(data_23),
        .data_24(data_24),
        .data_25(data_25),
        .data_26(data_26),
        .data_27(data_27),
        .data_28(data_28),
        .data_29(data_29),
        .data_30(data_30),
        .data_31(data_31),
        .data_32(data_32),
        .data_33(data_33),
        .sort_0(sort_0),
        .sort_1(sort_1),
        .sort_2(sort_2),
        .sort_3(sort_3),
        .sort_4(sort_4),
        .sort_5(sort_5),
        .sort_6(sort_6),
        .sort_7(sort_7),
        .sort_8(sort_8),
        .sort_9(sort_9),
        .sort_10(sort_10),
        .sort_11(sort_11),
        .sort_12(sort_12),
        .sort_13(sort_13),
        .sort_14(sort_14),
        .sort_15(sort_15),
        .sort_16(sort_16),
        .sort_17(sort_17),
        .sort_18(sort_18),
        .sort_19(sort_19),
        .sort_20(sort_20),
        .sort_21(sort_21),
        .sort_22(sort_22),
        .sort_23(sort_23),
        .sort_24(sort_24),
        .sort_25(sort_25),
        .sort_26(sort_26),
        .sort_27(sort_27),
        .sort_28(sort_28),
        .sort_29(sort_29),
        .sort_30(sort_30),
        .sort_31(sort_31),
        .sort_32(sort_32),
        .sort_33(sort_33)
    );

    // Apply random inputs
    initial begin
        repeat (100) begin
            @(posedge clk);
            data_0 = $urandom;
            data_1 = $urandom;
            data_2 = $urandom;
            data_3 = $urandom;
            data_4 = $urandom;
            data_5 = $urandom;
            data_6 = $urandom;
            data_7 = $urandom;
            data_8 = $urandom;
            data_9 = $urandom;
            data_10 = $urandom;
            data_11 = $urandom;
            data_12 = $urandom;
            data_13 = $urandom;
            data_14 = $urandom;
            data_15 = $urandom;
            data_16 = $urandom;
            data_17 = $urandom;
            data_18 = $urandom;
            data_19 = $urandom;
            data_20 = $urandom;
            data_21 = $urandom;
            data_22 = $urandom;
            data_23 = $urandom;
            data_24 = $urandom;
            data_25 = $urandom;
            data_26 = $urandom;
            data_27 = $urandom;
            data_28 = $urandom;
            data_29 = $urandom;
            data_30 = $urandom;
            data_31 = $urandom;
            data_32 = $urandom;
            data_33 = $urandom;
        end
        #100 $finish;
    end

    // Verification logic
    localparam int latency = 0;
    integer cycle_count = 0;
    integer success_count = 0;
    integer failure_count = 0;
    always @(posedge clk) begin
        cycle_count <= cycle_count + 1;
        if (cycle_count > latency) begin
            if (sort_0 <= sort_1 && sort_1 <= sort_2 && sort_2 <= sort_3 && sort_3 <= sort_4 && sort_4 <= sort_5 && sort_5 <= sort_6 && sort_6 <= sort_7 && sort_7 <= sort_8 && sort_8 <= sort_9 && sort_9 <= sort_10 && sort_10 <= sort_11 && sort_11 <= sort_12 && sort_12 <= sort_13 && sort_13 <= sort_14 && sort_14 <= sort_15 && sort_15 <= sort_16 && sort_16 <= sort_17 && sort_17 <= sort_18 && sort_18 <= sort_19 && sort_19 <= sort_20 && sort_20 <= sort_21 && sort_21 <= sort_22 && sort_22 <= sort_23 && sort_23 <= sort_24 && sort_24 <= sort_25 && sort_25 <= sort_26 && sort_26 <= sort_27 && sort_27 <= sort_28 && sort_28 <= sort_29 && sort_29 <= sort_30 && sort_30 <= sort_31 && sort_31 <= sort_32 && sort_32 <= sort_33) begin
                success_count <= success_count + 1;
            end else begin
                failure_count <= failure_count + 1;
            end
            $display("Cycle: %0d, Success: %0d, Failure: %0d", cycle_count, success_count, failure_count);
        end
    end

endmodule